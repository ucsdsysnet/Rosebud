module table_000000010(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b00010100001: match <= 1'b1;
      11'b010000010??: match <= 1'b1;
      11'b0010011????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_000000100(input clk, input rst, input [13:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      14'b01110101011000: match <= 1'b1;
      14'b01110101011001: match <= 1'b1;
      14'b0111000110000?: match <= 1'b1;
      14'b0111011110010?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_000001011(input clk, input rst, input [13:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      14'b01111000000101: match <= 1'b1;
      14'b0110100000001?: match <= 1'b1;
      14'b0110111001111?: match <= 1'b1;
      14'b0000110100????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_000110001(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b00010010001: match <= 1'b1;
      11'b01010101101: match <= 1'b1;
      11'b1101001000?: match <= 1'b1;
      11'b1101100000?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_000110110(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b11111101010: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_000110111(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0010010: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_000111110(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b000111001000001: match <= 1'b1;
      15'b0101000100111??: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001001000(input clk, input rst, input [11:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      12'b000000000001: match <= 1'b1;
      12'b01001010011?: match <= 1'b1;
      12'b1110100?????: match <= 1'b1;
      12'b1110111?????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001001011(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b001110010101101: match <= 1'b1;
      15'b00111000100000?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001010010(input clk, input rst, input [11:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      12'b100110111110: match <= 1'b1;
      12'b100100000???: match <= 1'b1;
      12'b10111011????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001010100(input clk, input rst, input [9:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      10'b0000000001: match <= 1'b1;
      10'b110000000?: match <= 1'b1;
      10'b00000011??: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001010101(input clk, input rst, input [2:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      3'b000: match <= 1'b1;
      3'b010: match <= 1'b1;
      3'b101: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001010111(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1100101001101: match <= 1'b1;
      13'b1111010011101: match <= 1'b1;
      13'b1111100010100: match <= 1'b1;
      13'b1101100??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001011010(input clk, input rst, input [13:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      14'b10100001111100: match <= 1'b1;
      14'b10100001111101: match <= 1'b1;
      14'b0000100100000?: match <= 1'b1;
      14'b0000100100010?: match <= 1'b1;
      14'b0000110001100?: match <= 1'b1;
      14'b0001001100101?: match <= 1'b1;
      14'b0001011101111?: match <= 1'b1;
      14'b1000001001000?: match <= 1'b1;
      14'b1000001011110?: match <= 1'b1;
      14'b1000001101111?: match <= 1'b1;
      14'b1000011111101?: match <= 1'b1;
      14'b1010000000111?: match <= 1'b1;
      14'b1010000010100?: match <= 1'b1;
      14'b1010110000101?: match <= 1'b1;
      14'b1110010111100?: match <= 1'b1;
      14'b1110111001010?: match <= 1'b1;
      14'b1111001110011?: match <= 1'b1;
      14'b01110110110???: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001011011(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0011111001110: match <= 1'b1;
      13'b101110001????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001011100(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b110011010110001: match <= 1'b1;
      15'b110011010111110: match <= 1'b1;
      15'b11001101011001?: match <= 1'b1;
      15'b11001101011011?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001011101(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0101110110011: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001100011(input clk, input rst, input [9:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      10'b0011100101: match <= 1'b1;
      10'b110111001?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001110100(input clk, input rst, input [5:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      6'b000111: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001110111(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0011001001111: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001111001(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b1101001: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001111010(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b010110111111011: match <= 1'b1;
      15'b0001011111?????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_001111110(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b110000111011011: match <= 1'b1;
      15'b10000100011110?: match <= 1'b1;
      15'b11000011101110?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010000000(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b00011110000: match <= 1'b1;
      11'b10001010001: match <= 1'b1;
      11'b10111001110: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010000001(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b11110101001: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010000010(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b11000010011: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010000011(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b100010011100101: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010000111(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b10101010111: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010001000(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b10000100011: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010001010(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b00010000100: match <= 1'b1;
      11'b00010000110: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010010000(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b00000011110: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010010100(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1110010100101: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010011001(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b01111110000: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010011010(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b010010000111110: match <= 1'b1;
      15'b101000101010110: match <= 1'b1;
      15'b101000101011001: match <= 1'b1;
      15'b10100010101010?: match <= 1'b1;
      15'b10100010101101?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010100111(input clk, input rst, input [8:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      9'b010111100: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010101000(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0100110000001: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010101001(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1101110101000: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010101010(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b111100100100111: match <= 1'b1;
      15'b1011100011111??: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010101011(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1010001000001: match <= 1'b1;
      13'b1010001010010: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010101100(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b110100000000010: match <= 1'b1;
      15'b110100100000010: match <= 1'b1;
      15'b110100100000110: match <= 1'b1;
      15'b110100110110000: match <= 1'b1;
      15'b110100110110010: match <= 1'b1;
      15'b110100110111010: match <= 1'b1;
      15'b110100111100101: match <= 1'b1;
      15'b110100111100110: match <= 1'b1;
      15'b110101000001010: match <= 1'b1;
      15'b110101000001101: match <= 1'b1;
      15'b110101001101001: match <= 1'b1;
      15'b110101001101101: match <= 1'b1;
      15'b110101001110110: match <= 1'b1;
      15'b110101101001000: match <= 1'b1;
      15'b110101111000001: match <= 1'b1;
      15'b01101110010100?: match <= 1'b1;
      15'b01101110010101?: match <= 1'b1;
      15'b11010000000000?: match <= 1'b1;
      15'b11010001101010?: match <= 1'b1;
      15'b11010001101111?: match <= 1'b1;
      15'b11010001110000?: match <= 1'b1;
      15'b11010011011100?: match <= 1'b1;
      15'b11010011111001?: match <= 1'b1;
      15'b11010100000111?: match <= 1'b1;
      15'b11010100101111?: match <= 1'b1;
      15'b11010100110101?: match <= 1'b1;
      15'b11010100110111?: match <= 1'b1;
      15'b11010100111001?: match <= 1'b1;
      15'b11010100111010?: match <= 1'b1;
      15'b11010101000101?: match <= 1'b1;
      15'b11010101000110?: match <= 1'b1;
      15'b11010101010111?: match <= 1'b1;
      15'b11010111100001?: match <= 1'b1;
      15'b0111110000111??: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010110001(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1011010001010: match <= 1'b1;
      13'b1011010100101: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010110010(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b010000000101011: match <= 1'b1;
      15'b010000010101010: match <= 1'b1;
      15'b010000011001010: match <= 1'b1;
      15'b010000101110100: match <= 1'b1;
      15'b010000110000110: match <= 1'b1;
      15'b010000111001110: match <= 1'b1;
      15'b010001000000000: match <= 1'b1;
      15'b010001000000100: match <= 1'b1;
      15'b010001001100110: match <= 1'b1;
      15'b010001100110110: match <= 1'b1;
      15'b010001101011001: match <= 1'b1;
      15'b010001101011010: match <= 1'b1;
      15'b010010010001000: match <= 1'b1;
      15'b010010010001101: match <= 1'b1;
      15'b010010101011110: match <= 1'b1;
      15'b010010101100000: match <= 1'b1;
      15'b010010110000001: match <= 1'b1;
      15'b010010110000110: match <= 1'b1;
      15'b010011011110000: match <= 1'b1;
      15'b010011101000101: match <= 1'b1;
      15'b010011111010100: match <= 1'b1;
      15'b010011111010111: match <= 1'b1;
      15'b010011111110001: match <= 1'b1;
      15'b010100010001010: match <= 1'b1;
      15'b010100011001111: match <= 1'b1;
      15'b010100011010001: match <= 1'b1;
      15'b010100100011011: match <= 1'b1;
      15'b010100100110001: match <= 1'b1;
      15'b010100110111101: match <= 1'b1;
      15'b010101000001010: match <= 1'b1;
      15'b010101010011010: match <= 1'b1;
      15'b010110101010010: match <= 1'b1;
      15'b010111000101111: match <= 1'b1;
      15'b01000010010111?: match <= 1'b1;
      15'b01000011100011?: match <= 1'b1;
      15'b01000011100100?: match <= 1'b1;
      15'b01000011111101?: match <= 1'b1;
      15'b01000011111111?: match <= 1'b1;
      15'b01000100110100?: match <= 1'b1;
      15'b01001000010011?: match <= 1'b1;
      15'b01001001000101?: match <= 1'b1;
      15'b01001010101110?: match <= 1'b1;
      15'b01001011000001?: match <= 1'b1;
      15'b01001011000010?: match <= 1'b1;
      15'b01010001000110?: match <= 1'b1;
      15'b01010010001110?: match <= 1'b1;
      15'b01010010011001?: match <= 1'b1;
      15'b01010011011111?: match <= 1'b1;
      15'b01010101001100?: match <= 1'b1;
      15'b0101110000010??: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010110111(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b100100010000101: match <= 1'b1;
      15'b101110010100011: match <= 1'b1;
      15'b110100000010010: match <= 1'b1;
      15'b111011011001000: match <= 1'b1;
      15'b11010111000001?: match <= 1'b1;
      15'b0000100101001??: match <= 1'b1;
      15'b1000101110001??: match <= 1'b1;
      15'b1001000000011??: match <= 1'b1;
      15'b1001000111110??: match <= 1'b1;
      15'b1011010111011??: match <= 1'b1;
      15'b1100101001101??: match <= 1'b1;
      15'b1110011101100??: match <= 1'b1;
      15'b111011010110???: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010111000(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1110110010100: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010111010(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b111001000110011: match <= 1'b1;
      15'b111001000110110: match <= 1'b1;
      15'b111001100111011: match <= 1'b1;
      15'b111100000100010: match <= 1'b1;
      15'b111100000101110: match <= 1'b1;
      15'b11100100011010?: match <= 1'b1;
      15'b11100100011101?: match <= 1'b1;
      15'b11101110111011?: match <= 1'b1;
      15'b11101110111100?: match <= 1'b1;
      15'b11101110111110?: match <= 1'b1;
      15'b1110010001111??: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_010111101(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0000011111001: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011000000(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b01011011001: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011001010(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0101010: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011001011(input clk, input rst, input [9:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      10'b1001011100: match <= 1'b1;
      10'b000011????: match <= 1'b1;
      10'b111100????: match <= 1'b1;
      10'b10000?????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011001101(input clk, input rst, input [9:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      10'b1000100011: match <= 1'b1;
      10'b1010011111: match <= 1'b1;
      10'b1010100111: match <= 1'b1;
      10'b1100100???: match <= 1'b1;
      10'b1101000???: match <= 1'b1;
      10'b1110000???: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011001110(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0001110110100: match <= 1'b1;
      13'b0010111000010: match <= 1'b1;
      13'b0010111011111: match <= 1'b1;
      13'b0011110000011: match <= 1'b1;
      13'b0100000100001: match <= 1'b1;
      13'b0100100010000: match <= 1'b1;
      13'b0111011010111: match <= 1'b1;
      13'b1001001101011: match <= 1'b1;
      13'b1001011001001: match <= 1'b1;
      13'b1001100011000: match <= 1'b1;
      13'b1001100100000: match <= 1'b1;
      13'b1001101001000: match <= 1'b1;
      13'b1100011000000: match <= 1'b1;
      13'b1100100101010: match <= 1'b1;
      13'b0100000??????: match <= 1'b1;
      13'b0100010??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011001111(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b000011110010000: match <= 1'b1;
      15'b00001101001000?: match <= 1'b1;
      15'b1000101111100??: match <= 1'b1;
      15'b1000111010110??: match <= 1'b1;
      15'b1010010111101??: match <= 1'b1;
      15'b1010111010100??: match <= 1'b1;
      15'b1100001010010??: match <= 1'b1;
      15'b1100001100000??: match <= 1'b1;
      15'b1100010110000??: match <= 1'b1;
      15'b1100100001111??: match <= 1'b1;
      15'b1100101001001??: match <= 1'b1;
      15'b1100110100100??: match <= 1'b1;
      15'b1101000100010??: match <= 1'b1;
      15'b1101000101011??: match <= 1'b1;
      15'b1101100001000??: match <= 1'b1;
      15'b1101111001110??: match <= 1'b1;
      15'b1110011000010??: match <= 1'b1;
      15'b0101011111?????: match <= 1'b1;
      15'b0101110111?????: match <= 1'b1;
      15'b0110100111?????: match <= 1'b1;
      15'b0111101111?????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011010001(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b101101011101111: match <= 1'b1;
      15'b0011001111101??: match <= 1'b1;
      15'b00011110001????: match <= 1'b1;
      15'b11100111100????: match <= 1'b1;
      15'b1001111010?????: match <= 1'b1;
      15'b1111010110?????: match <= 1'b1;
      15'b110100100??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011010100(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b1011111: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011010111(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b01101100111: match <= 1'b1;
      11'b01101101111: match <= 1'b1;
      11'b01111101010: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011011100(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0101001: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011011111(input clk, input rst, input [9:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      10'b1011111110: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011100011(input clk, input rst, input [9:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      10'b1010100100: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011101001(input clk, input rst, input [5:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      6'b001000: match <= 1'b1;
      6'b001001: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011101010(input clk, input rst, input [7:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      8'b01110100: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011101110(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0111010: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011101111(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b1101000: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011110000(input clk, input rst, input [5:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      6'b011000: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011110100(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0001000: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011110101(input clk, input rst, input [8:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      9'b000000100: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011110111(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b00010000101: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011111000(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0010100: match <= 1'b1;
      7'b100010?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011111001(input clk, input rst, input [8:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      9'b001110100: match <= 1'b1;
      9'b1110010??: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011111010(input clk, input rst, input [8:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      9'b001111111: match <= 1'b1;
      9'b011101000: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_011111011(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0101001: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100000000(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0011000: match <= 1'b1;
      7'b1010101: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100000100(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0010101: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100000101(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0010100: match <= 1'b1;
      7'b1000100: match <= 1'b1;
      7'b1011110: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100000110(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1101100000100: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100000111(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0001111: match <= 1'b1;
      7'b1001000: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100001001(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1111111100001: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100001100(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0010010: match <= 1'b1;
      7'b0010110: match <= 1'b1;
      7'b0010111: match <= 1'b1;
      7'b0100001: match <= 1'b1;
      7'b1111111: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100001101(input clk, input rst, input [8:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      9'b010110011: match <= 1'b1;
      9'b0101100??: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100010010(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0010011: match <= 1'b1;
      7'b0011111: match <= 1'b1;
      7'b0100001: match <= 1'b1;
      7'b0110111: match <= 1'b1;
      7'b1001000: match <= 1'b1;
      7'b1001100: match <= 1'b1;
      7'b1101001: match <= 1'b1;
      7'b1110010: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100010011(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0101011: match <= 1'b1;
      7'b1011010: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100010100(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0100100010111: match <= 1'b1;
      13'b0100100100010: match <= 1'b1;
      13'b0111011000001: match <= 1'b1;
      13'b0111011110011: match <= 1'b1;
      13'b1011110100100: match <= 1'b1;
      13'b1011110110110: match <= 1'b1;
      13'b1100001100111: match <= 1'b1;
      13'b1111010110000: match <= 1'b1;
      13'b0011111??????: match <= 1'b1;
      13'b0110100??????: match <= 1'b1;
      13'b1111101??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100010101(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0111001011101: match <= 1'b1;
      13'b0111010110100: match <= 1'b1;
      13'b1011011101011: match <= 1'b1;
      13'b1011000??????: match <= 1'b1;
      13'b1111001??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100010110(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0101100: match <= 1'b1;
      7'b1010001: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100010111(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0111100: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100011000(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b10100100110: match <= 1'b1;
      11'b1010010010?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100011001(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0100111: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100011010(input clk, input rst, input [13:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      14'b11000100100010: match <= 1'b1;
      14'b11000100100011: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100011011(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b10011101000: match <= 1'b1;
      11'b0110010????: match <= 1'b1;
      11'b1111101????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100011100(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b1100110: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100011110(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0000000111011: match <= 1'b1;
      13'b0110001??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100011111(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0000111: match <= 1'b1;
      7'b0001000: match <= 1'b1;
      7'b1111101: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100100011(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b1100111: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100100100(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0000011: match <= 1'b1;
      7'b0110011: match <= 1'b1;
      7'b1101010: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100100101(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0110111: match <= 1'b1;
      7'b1001010: match <= 1'b1;
      7'b1111100: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100100110(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1001110111000: match <= 1'b1;
      13'b0000111??????: match <= 1'b1;
      13'b1110111??????: match <= 1'b1;
      13'b00100????????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100101001(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0010100: match <= 1'b1;
      7'b0011010: match <= 1'b1;
      7'b0110010: match <= 1'b1;
      7'b0111001: match <= 1'b1;
      7'b1111000: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100101010(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b1110110: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100101011(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b1001111: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100101100(input clk, input rst, input [7:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      8'b00101101: match <= 1'b1;
      8'b0001010?: match <= 1'b1;
      8'b0011001?: match <= 1'b1;
      8'b0101000?: match <= 1'b1;
      8'b1111001?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100101101(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0000001110101: match <= 1'b1;
      13'b0000001111001: match <= 1'b1;
      13'b1110010011110: match <= 1'b1;
      13'b1110010100100: match <= 1'b1;
      13'b0001101??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100101111(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b1010100: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100110000(input clk, input rst, input [13:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      14'b10110011110010: match <= 1'b1;
      14'b10110011110011: match <= 1'b1;
      14'b1101101???????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100110001(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0010011: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100110010(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0001110: match <= 1'b1;
      7'b1011101: match <= 1'b1;
      7'b01101??: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100110110(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0101000: match <= 1'b1;
      7'b1000010: match <= 1'b1;
      7'b1000111: match <= 1'b1;
      7'b1001001: match <= 1'b1;
      7'b1101100: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100110111(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0011111: match <= 1'b1;
      7'b1101001: match <= 1'b1;
      7'b1101011: match <= 1'b1;
      7'b1111001: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100111000(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b1100000: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100111001(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1100101100001: match <= 1'b1;
      13'b110010110001?: match <= 1'b1;
      13'b110100110000?: match <= 1'b1;
      13'b110100110001?: match <= 1'b1;
      13'b11001011001??: match <= 1'b1;
      13'b11010011001??: match <= 1'b1;
      13'b1100101101???: match <= 1'b1;
      13'b1101001101???: match <= 1'b1;
      13'b1101001110???: match <= 1'b1;
      13'b1101001111???: match <= 1'b1;
      13'b110010111????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100111010(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b1110011: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100111011(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0100010: match <= 1'b1;
      7'b0111010: match <= 1'b1;
      7'b1000011: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100111100(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0110110: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100111101(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b1111001: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100111110(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b1010000: match <= 1'b1;
      7'b1010101: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_100111111(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0101110: match <= 1'b1;
      7'b1011011: match <= 1'b1;
      7'b1100101: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101000000(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0001110: match <= 1'b1;
      7'b0010101: match <= 1'b1;
      7'b1110011: match <= 1'b1;
      7'b1110100: match <= 1'b1;
      7'b1110101: match <= 1'b1;
      7'b1111001: match <= 1'b1;
      7'b1111010: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101000001(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0110100: match <= 1'b1;
      7'b0110101: match <= 1'b1;
      7'b0111000: match <= 1'b1;
      7'b0111100: match <= 1'b1;
      7'b1001000: match <= 1'b1;
      7'b1101011: match <= 1'b1;
      7'b1110000: match <= 1'b1;
      7'b1111111: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101000010(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0000000010001: match <= 1'b1;
      13'b0000000000???: match <= 1'b1;
      13'b0000001??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101000101(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1010000011111: match <= 1'b1;
      13'b1010100101111: match <= 1'b1;
      13'b1111001000101: match <= 1'b1;
      13'b1111011010111: match <= 1'b1;
      13'b101111010000?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101000110(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b010111100010011: match <= 1'b1;
      15'b011010111110111: match <= 1'b1;
      15'b1111111111?????: match <= 1'b1;
      15'b0110010????????: match <= 1'b1;
      15'b0111011????????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101000111(input clk, input rst, input [9:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      10'b0000000111: match <= 1'b1;
      10'b1011000000: match <= 1'b1;
      10'b1000101???: match <= 1'b1;
      10'b1000110???: match <= 1'b1;
      10'b1111010???: match <= 1'b1;
      10'b1111110???: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101001000(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0000110: match <= 1'b1;
      7'b1001111: match <= 1'b1;
      7'b1011000: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101001001(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0001001: match <= 1'b1;
      7'b0011011: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101001010(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0000011: match <= 1'b1;
      7'b0011001: match <= 1'b1;
      7'b1100110: match <= 1'b1;
      7'b01101??: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101001011(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b1001101: match <= 1'b1;
      7'b1010001: match <= 1'b1;
      7'b1100111: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101001100(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b1011101: match <= 1'b1;
      7'b1110101: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101001110(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b10100101001: match <= 1'b1;
      11'b100101000??: match <= 1'b1;
      11'b1100111????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101001111(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1111001110010: match <= 1'b1;
      13'b110000000110?: match <= 1'b1;
      13'b11000000010??: match <= 1'b1;
      13'b0100000011???: match <= 1'b1;
      13'b1100000000???: match <= 1'b1;
      13'b0011110??????: match <= 1'b1;
      13'b0100010??????: match <= 1'b1;
      13'b0101111??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101010000(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0000000110101: match <= 1'b1;
      13'b1011010011000: match <= 1'b1;
      13'b1000000??????: match <= 1'b1;
      13'b1001100??????: match <= 1'b1;
      13'b101000???????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101010001(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b001011100000110: match <= 1'b1;
      15'b001011100101011: match <= 1'b1;
      15'b001011100110110: match <= 1'b1;
      15'b001011110010001: match <= 1'b1;
      15'b001011110011101: match <= 1'b1;
      15'b001011111111110: match <= 1'b1;
      15'b00101110000010?: match <= 1'b1;
      15'b00101110011010?: match <= 1'b1;
      15'b00101110100010?: match <= 1'b1;
      15'b00101111001001?: match <= 1'b1;
      15'b00101111001111?: match <= 1'b1;
      15'b00101111101110?: match <= 1'b1;
      15'b0010111000000??: match <= 1'b1;
      15'b0010111001011??: match <= 1'b1;
      15'b0010111001100??: match <= 1'b1;
      15'b0010111010000??: match <= 1'b1;
      15'b0010111100101??: match <= 1'b1;
      15'b0010111100110??: match <= 1'b1;
      15'b0010111101110??: match <= 1'b1;
      15'b0010111110110??: match <= 1'b1;
      15'b0010111111110??: match <= 1'b1;
      15'b0110101001101??: match <= 1'b1;
      15'b1000011010011??: match <= 1'b1;
      15'b1000100111011??: match <= 1'b1;
      15'b1000100111100??: match <= 1'b1;
      15'b1001101010010??: match <= 1'b1;
      15'b1100011100000??: match <= 1'b1;
      15'b1100011100011??: match <= 1'b1;
      15'b001011100100???: match <= 1'b1;
      15'b001011100111???: match <= 1'b1;
      15'b001011101001???: match <= 1'b1;
      15'b001011110110???: match <= 1'b1;
      15'b001011111010???: match <= 1'b1;
      15'b001011111101???: match <= 1'b1;
      15'b001011111110???: match <= 1'b1;
      15'b00101110101????: match <= 1'b1;
      15'b00101111000????: match <= 1'b1;
      15'b00101111010????: match <= 1'b1;
      15'b00101111100????: match <= 1'b1;
      15'b0010111011?????: match <= 1'b1;
      15'b0000001????????: match <= 1'b1;
      15'b1000110????????: match <= 1'b1;
      15'b1001110????????: match <= 1'b1;
      15'b1010011????????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101010011(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1101111100110: match <= 1'b1;
      13'b0001000111???: match <= 1'b1;
      13'b0000001??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101010100(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1010011111010: match <= 1'b1;
      13'b1000011??????: match <= 1'b1;
      13'b1110001??????: match <= 1'b1;
      13'b1111000??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101010101(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1110100001010: match <= 1'b1;
      13'b1110100111100: match <= 1'b1;
      13'b1110111110111: match <= 1'b1;
      13'b0110011??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101010110(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0011010: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101011110(input clk, input rst, input [8:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      9'b110011101: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101100000(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b110111110101110: match <= 1'b1;
      15'b111100100001110: match <= 1'b1;
      15'b111111011000010: match <= 1'b1;
      15'b11111101100000?: match <= 1'b1;
      15'b1110100111010??: match <= 1'b1;
      15'b110000001011???: match <= 1'b1;
      15'b110011001111???: match <= 1'b1;
      15'b110011111110???: match <= 1'b1;
      15'b0111000110?????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101100001(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b101111101110110: match <= 1'b1;
      15'b10111110111010?: match <= 1'b1;
      15'b10111111010000?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101100011(input clk, input rst, input [11:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      12'b110101010001: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101100101(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1010101101100: match <= 1'b1;
      13'b101010010111?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101100110(input clk, input rst, input [7:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      8'b01111110: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101101001(input clk, input rst, input [8:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      9'b011001011: match <= 1'b1;
      9'b11011????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101101011(input clk, input rst, input [11:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      12'b110000011000: match <= 1'b1;
      12'b110000011011: match <= 1'b1;
      12'b110100110011: match <= 1'b1;
      12'b01011101101?: match <= 1'b1;
      12'b01011101110?: match <= 1'b1;
      12'b01011101111?: match <= 1'b1;
      12'b11010011000?: match <= 1'b1;
      12'b1100000000??: match <= 1'b1;
      12'b1100000001??: match <= 1'b1;
      12'b1100000010??: match <= 1'b1;
      12'b1101001101??: match <= 1'b1;
      12'b011000101???: match <= 1'b1;
      12'b011110100???: match <= 1'b1;
      12'b110100010???: match <= 1'b1;
      12'b110100011???: match <= 1'b1;
      12'b110100100???: match <= 1'b1;
      12'b110100101???: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101110010(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b011110011001001: match <= 1'b1;
      15'b011111100100011: match <= 1'b1;
      15'b100000000010111: match <= 1'b1;
      15'b100110111111000: match <= 1'b1;
      15'b111010010101111: match <= 1'b1;
      15'b01111001100101?: match <= 1'b1;
      15'b11101001010110?: match <= 1'b1;
      15'b0010101000010??: match <= 1'b1;
      15'b0011110101010??: match <= 1'b1;
      15'b0110111000001??: match <= 1'b1;
      15'b0110111100011??: match <= 1'b1;
      15'b1010000011100??: match <= 1'b1;
      15'b1010001101101??: match <= 1'b1;
      15'b1100110001100??: match <= 1'b1;
      15'b1101001001110??: match <= 1'b1;
      15'b1101110000000??: match <= 1'b1;
      15'b1111000000010??: match <= 1'b1;
      15'b1111010100000??: match <= 1'b1;
      15'b1111100000000??: match <= 1'b1;
      15'b1111111001011??: match <= 1'b1;
      15'b1111111001110??: match <= 1'b1;
      15'b1111111010001??: match <= 1'b1;
      15'b1111111010011??: match <= 1'b1;
      15'b111101111111???: match <= 1'b1;
      15'b111110000111???: match <= 1'b1;
      15'b111111010100???: match <= 1'b1;
      15'b0000000011?????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101110011(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b100000101011010: match <= 1'b1;
      15'b101011101110001: match <= 1'b1;
      15'b11011011110001?: match <= 1'b1;
      15'b0000001000010??: match <= 1'b1;
      15'b0000001110100??: match <= 1'b1;
      15'b0000010001001??: match <= 1'b1;
      15'b0000100000010??: match <= 1'b1;
      15'b0000110001100??: match <= 1'b1;
      15'b0010000101101??: match <= 1'b1;
      15'b0010011100011??: match <= 1'b1;
      15'b0011100010111??: match <= 1'b1;
      15'b0100001100101??: match <= 1'b1;
      15'b0100101000110??: match <= 1'b1;
      15'b0110100110000??: match <= 1'b1;
      15'b0111000110000??: match <= 1'b1;
      15'b0111001001100??: match <= 1'b1;
      15'b1000010011001??: match <= 1'b1;
      15'b1010111100001??: match <= 1'b1;
      15'b1100011110010??: match <= 1'b1;
      15'b1100110001011??: match <= 1'b1;
      15'b1101010010000??: match <= 1'b1;
      15'b1101100111010??: match <= 1'b1;
      15'b1101101011010??: match <= 1'b1;
      15'b1101101110111??: match <= 1'b1;
      15'b1101110101100??: match <= 1'b1;
      15'b1111000100001??: match <= 1'b1;
      15'b001110001011???: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101110100(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b10000010111: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101110101(input clk, input rst, input [8:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      9'b011001100: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101111001(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b101000001101101: match <= 1'b1;
      15'b101010011111110: match <= 1'b1;
      15'b101010100010111: match <= 1'b1;
      15'b101011001011110: match <= 1'b1;
      15'b101011001011111: match <= 1'b1;
      15'b101011010001100: match <= 1'b1;
      15'b101011010011011: match <= 1'b1;
      15'b101011011000001: match <= 1'b1;
      15'b111000111010011: match <= 1'b1;
      15'b111011111100110: match <= 1'b1;
      15'b10101011100111?: match <= 1'b1;
      15'b10101011101011?: match <= 1'b1;
      15'b1010000001100??: match <= 1'b1;
      15'b1010000001101??: match <= 1'b1;
      15'b1010000110111??: match <= 1'b1;
      15'b1010101111110??: match <= 1'b1;
      15'b1010101111111??: match <= 1'b1;
      15'b101000101111???: match <= 1'b1;
      15'b0101100101?????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101111100(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1100111101111: match <= 1'b1;
      13'b11001100010??: match <= 1'b1;
      13'b11110111101??: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_101111101(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0111001011000: match <= 1'b1;
      13'b0111001011011: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110000000(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b000010101100111: match <= 1'b1;
      15'b000110010000011: match <= 1'b1;
      15'b001101000011001: match <= 1'b1;
      15'b010100000011101: match <= 1'b1;
      15'b010101110100000: match <= 1'b1;
      15'b010101110101111: match <= 1'b1;
      15'b010101110111000: match <= 1'b1;
      15'b011011001101110: match <= 1'b1;
      15'b100001100010000: match <= 1'b1;
      15'b110000010010010: match <= 1'b1;
      15'b110010100101100: match <= 1'b1;
      15'b110010110110101: match <= 1'b1;
      15'b00111111101010?: match <= 1'b1;
      15'b11001011111100?: match <= 1'b1;
      15'b010101110110???: match <= 1'b1;
      15'b110010111001???: match <= 1'b1;
      15'b110010111110???: match <= 1'b1;
      15'b11001011101????: match <= 1'b1;
      15'b11001011110????: match <= 1'b1;
      15'b0010110????????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110000001(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b000010100000011: match <= 1'b1;
      15'b001100011000010: match <= 1'b1;
      15'b001101000001011: match <= 1'b1;
      15'b010000000101100: match <= 1'b1;
      15'b011111000110001: match <= 1'b1;
      15'b011111001100001: match <= 1'b1;
      15'b100001110010110: match <= 1'b1;
      15'b100010101010111: match <= 1'b1;
      15'b100101111111100: match <= 1'b1;
      15'b100111001110010: match <= 1'b1;
      15'b110011101000010: match <= 1'b1;
      15'b110101010011100: match <= 1'b1;
      15'b110101010111101: match <= 1'b1;
      15'b111010101100101: match <= 1'b1;
      15'b111010110111100: match <= 1'b1;
      15'b111010111111000: match <= 1'b1;
      15'b111101111100111: match <= 1'b1;
      15'b101101101111???: match <= 1'b1;
      15'b101101111010???: match <= 1'b1;
      15'b10110111100????: match <= 1'b1;
      15'b11000100001????: match <= 1'b1;
      15'b11111000001????: match <= 1'b1;
      15'b1100101001?????: match <= 1'b1;
      15'b101101110??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110000010(input clk, input rst, input [13:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      14'b00111101111111: match <= 1'b1;
      14'b01000000100001: match <= 1'b1;
      14'b0101110101011?: match <= 1'b1;
      14'b00110010011???: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110000011(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b110010001011011: match <= 1'b1;
      15'b0010111101000??: match <= 1'b1;
      15'b11111100011????: match <= 1'b1;
      15'b11100110???????: match <= 1'b1;
      15'b0001011????????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110000100(input clk, input rst, input [13:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      14'b00001010101111: match <= 1'b1;
      14'b01010010011110: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110000101(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b001001110001100: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110000111(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b011011000111001: match <= 1'b1;
      15'b1010010011?????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110001000(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b000000101101101: match <= 1'b1;
      15'b000101000111101: match <= 1'b1;
      15'b00010100011111?: match <= 1'b1;
      15'b01111011100????: match <= 1'b1;
      15'b0001010010?????: match <= 1'b1;
      15'b000111101??????: match <= 1'b1;
      15'b01010101???????: match <= 1'b1;
      15'b0111110????????: match <= 1'b1;
      15'b0111111????????: match <= 1'b1;
      15'b00100??????????: match <= 1'b1;
      15'b01101??????????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110001001(input clk, input rst, input [8:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      9'b100000011: match <= 1'b1;
      9'b100111101: match <= 1'b1;
      9'b1000001??: match <= 1'b1;
      9'b1110110??: match <= 1'b1;
      9'b100001???: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110001011(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1100111110100: match <= 1'b1;
      13'b0011010??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110001100(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b011011011101000: match <= 1'b1;
      15'b011111001000110: match <= 1'b1;
      15'b011111001001100: match <= 1'b1;
      15'b110001101110101: match <= 1'b1;
      15'b110011011011110: match <= 1'b1;
      15'b00011010000????: match <= 1'b1;
      15'b00011100000????: match <= 1'b1;
      15'b00101000001????: match <= 1'b1;
      15'b01011010010????: match <= 1'b1;
      15'b01110010100????: match <= 1'b1;
      15'b11000001110????: match <= 1'b1;
      15'b0101101010?????: match <= 1'b1;
      15'b011100001??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110001101(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b000010101111000: match <= 1'b1;
      15'b001010011010100: match <= 1'b1;
      15'b010000011001101: match <= 1'b1;
      15'b010100111001001: match <= 1'b1;
      15'b011000110101111: match <= 1'b1;
      15'b011000110110100: match <= 1'b1;
      15'b011000111010110: match <= 1'b1;
      15'b011001100010110: match <= 1'b1;
      15'b011100011000001: match <= 1'b1;
      15'b011100011010000: match <= 1'b1;
      15'b011101000011001: match <= 1'b1;
      15'b011101111000000: match <= 1'b1;
      15'b011111010101101: match <= 1'b1;
      15'b100011111010100: match <= 1'b1;
      15'b100101011101101: match <= 1'b1;
      15'b100111010001100: match <= 1'b1;
      15'b101010010000100: match <= 1'b1;
      15'b10010000000100?: match <= 1'b1;
      15'b0010111100110??: match <= 1'b1;
      15'b0110001101100??: match <= 1'b1;
      15'b100100000000???: match <= 1'b1;
      15'b100110000000???: match <= 1'b1;
      15'b00101110001????: match <= 1'b1;
      15'b01101010110????: match <= 1'b1;
      15'b0110010010?????: match <= 1'b1;
      15'b0110111001?????: match <= 1'b1;
      15'b001011101??????: match <= 1'b1;
      15'b011101101??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110001110(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b000010010010111: match <= 1'b1;
      15'b000010111000010: match <= 1'b1;
      15'b000010111100101: match <= 1'b1;
      15'b001101010001001: match <= 1'b1;
      15'b001101010110101: match <= 1'b1;
      15'b001101011001101: match <= 1'b1;
      15'b001101011001111: match <= 1'b1;
      15'b001101011111011: match <= 1'b1;
      15'b010000111011110: match <= 1'b1;
      15'b011110001100110: match <= 1'b1;
      15'b100011110001011: match <= 1'b1;
      15'b101010000110111: match <= 1'b1;
      15'b101010000111100: match <= 1'b1;
      15'b101100111000110: match <= 1'b1;
      15'b111100010100011: match <= 1'b1;
      15'b00001001110001?: match <= 1'b1;
      15'b00001001110010?: match <= 1'b1;
      15'b00001011001100?: match <= 1'b1;
      15'b1010100001110??: match <= 1'b1;
      15'b010011000000???: match <= 1'b1;
      15'b10001111100????: match <= 1'b1;
      15'b10010010100????: match <= 1'b1;
      15'b10101000001????: match <= 1'b1;
      15'b10110010001????: match <= 1'b1;
      15'b0011011001?????: match <= 1'b1;
      15'b1010100010?????: match <= 1'b1;
      15'b010001010??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110001111(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b010010010001000: match <= 1'b1;
      15'b010010111101101: match <= 1'b1;
      15'b010010111101110: match <= 1'b1;
      15'b010011011010001: match <= 1'b1;
      15'b011100001010010: match <= 1'b1;
      15'b011100011011111: match <= 1'b1;
      15'b100100111010100: match <= 1'b1;
      15'b110100101001110: match <= 1'b1;
      15'b110100101010101: match <= 1'b1;
      15'b110100101100000: match <= 1'b1;
      15'b110100101100101: match <= 1'b1;
      15'b111010101111011: match <= 1'b1;
      15'b111010110001010: match <= 1'b1;
      15'b111011000100011: match <= 1'b1;
      15'b111011010001001: match <= 1'b1;
      15'b111011011010101: match <= 1'b1;
      15'b111011011010111: match <= 1'b1;
      15'b111011011100010: match <= 1'b1;
      15'b111100011111110: match <= 1'b1;
      15'b01001101101011?: match <= 1'b1;
      15'b10001101011100?: match <= 1'b1;
      15'b0100110110010??: match <= 1'b1;
      15'b1000110101111??: match <= 1'b1;
      15'b100011010110???: match <= 1'b1;
      15'b110011001100???: match <= 1'b1;
      15'b111000100000???: match <= 1'b1;
      15'b111010000111???: match <= 1'b1;
      15'b111110100110???: match <= 1'b1;
      15'b01110011001????: match <= 1'b1;
      15'b10001101010????: match <= 1'b1;
      15'b10101000110????: match <= 1'b1;
      15'b10111110000????: match <= 1'b1;
      15'b11111010010????: match <= 1'b1;
      15'b11111011110????: match <= 1'b1;
      15'b11111100010????: match <= 1'b1;
      15'b0100101001?????: match <= 1'b1;
      15'b1000100110?????: match <= 1'b1;
      15'b1001000010?????: match <= 1'b1;
      15'b1100110010?????: match <= 1'b1;
      15'b1110001010?????: match <= 1'b1;
      15'b1111001010?????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110010000(input clk, input rst, input [13:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      14'b00000000011110: match <= 1'b1;
      14'b1000111011111?: match <= 1'b1;
      14'b011001011100??: match <= 1'b1;
      14'b0010110???????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110010001(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0111101001011: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110010011(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0010100101010: match <= 1'b1;
      13'b0101001??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110010100(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b001101101100010: match <= 1'b1;
      15'b001101101100011: match <= 1'b1;
      15'b001101110100001: match <= 1'b1;
      15'b001101110101000: match <= 1'b1;
      15'b00110110110000?: match <= 1'b1;
      15'b00110111010001?: match <= 1'b1;
      15'b0011011011001??: match <= 1'b1;
      15'b0011011011110??: match <= 1'b1;
      15'b0011011101001??: match <= 1'b1;
      15'b1010110000000??: match <= 1'b1;
      15'b0010100001?????: match <= 1'b1;
      15'b0010101010?????: match <= 1'b1;
      15'b0101000001?????: match <= 1'b1;
      15'b000000011??????: match <= 1'b1;
      15'b010100001??????: match <= 1'b1;
      15'b100010000??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110010101(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b00101000010: match <= 1'b1;
      11'b00101001011: match <= 1'b1;
      11'b01111010101: match <= 1'b1;
      11'b0110111000?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110010110(input clk, input rst, input [13:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      14'b00111110101100: match <= 1'b1;
      14'b01000100100011: match <= 1'b1;
      14'b0000010110010?: match <= 1'b1;
      14'b1010110111111?: match <= 1'b1;
      14'b0001001000????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110010111(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0101001000000: match <= 1'b1;
      13'b011111101????: match <= 1'b1;
      13'b100001100????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110011000(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b001101110011011: match <= 1'b1;
      15'b011010010111000: match <= 1'b1;
      15'b011010011111111: match <= 1'b1;
      15'b011111010110001: match <= 1'b1;
      15'b100101110010011: match <= 1'b1;
      15'b100101111100100: match <= 1'b1;
      15'b101000010100100: match <= 1'b1;
      15'b101000010110100: match <= 1'b1;
      15'b101000011000110: match <= 1'b1;
      15'b101011110001000: match <= 1'b1;
      15'b101011110101111: match <= 1'b1;
      15'b101011111000111: match <= 1'b1;
      15'b101011111101001: match <= 1'b1;
      15'b101100111100000: match <= 1'b1;
      15'b110101110000100: match <= 1'b1;
      15'b110101111010000: match <= 1'b1;
      15'b110101111101101: match <= 1'b1;
      15'b00100110010011?: match <= 1'b1;
      15'b11111101111010?: match <= 1'b1;
      15'b0001110010100??: match <= 1'b1;
      15'b101101110001???: match <= 1'b1;
      15'b111001110000???: match <= 1'b1;
      15'b01011000010????: match <= 1'b1;
      15'b01011001101????: match <= 1'b1;
      15'b01011001110????: match <= 1'b1;
      15'b01110010001????: match <= 1'b1;
      15'b10101100001????: match <= 1'b1;
      15'b10110001010????: match <= 1'b1;
      15'b11011101001????: match <= 1'b1;
      15'b11111100010????: match <= 1'b1;
      15'b0110100011?????: match <= 1'b1;
      15'b1101010110?????: match <= 1'b1;
      15'b110101010??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110011001(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b000000010010111: match <= 1'b1;
      15'b000000010110100: match <= 1'b1;
      15'b000001010100111: match <= 1'b1;
      15'b000001011000011: match <= 1'b1;
      15'b110000110011111: match <= 1'b1;
      15'b110000111010010: match <= 1'b1;
      15'b110111000100011: match <= 1'b1;
      15'b110111000101000: match <= 1'b1;
      15'b110111010001001: match <= 1'b1;
      15'b110111010101010: match <= 1'b1;
      15'b110111010110111: match <= 1'b1;
      15'b001001101000???: match <= 1'b1;
      15'b100001001000???: match <= 1'b1;
      15'b00000000010????: match <= 1'b1;
      15'b00000100001????: match <= 1'b1;
      15'b00100110110????: match <= 1'b1;
      15'b00100111111????: match <= 1'b1;
      15'b00111001100????: match <= 1'b1;
      15'b11010110001????: match <= 1'b1;
      15'b1111111001?????: match <= 1'b1;
      15'b110100000??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110011011(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b001011100111010: match <= 1'b1;
      15'b001011111011000: match <= 1'b1;
      15'b001111100101101: match <= 1'b1;
      15'b001111110101110: match <= 1'b1;
      15'b001111110110100: match <= 1'b1;
      15'b001111111001001: match <= 1'b1;
      15'b001111111110001: match <= 1'b1;
      15'b010011000101101: match <= 1'b1;
      15'b010011001001101: match <= 1'b1;
      15'b010011001010100: match <= 1'b1;
      15'b010011001010111: match <= 1'b1;
      15'b010011010000010: match <= 1'b1;
      15'b010011010101000: match <= 1'b1;
      15'b010011010110111: match <= 1'b1;
      15'b010011011010011: match <= 1'b1;
      15'b011110101000111: match <= 1'b1;
      15'b011110111001111: match <= 1'b1;
      15'b100111110000110: match <= 1'b1;
      15'b101001000011101: match <= 1'b1;
      15'b101001001101011: match <= 1'b1;
      15'b101001010001011: match <= 1'b1;
      15'b101001010101011: match <= 1'b1;
      15'b101001011111001: match <= 1'b1;
      15'b101001110101100: match <= 1'b1;
      15'b101001110110011: match <= 1'b1;
      15'b110100100010011: match <= 1'b1;
      15'b110100110011100: match <= 1'b1;
      15'b110100111011100: match <= 1'b1;
      15'b110110000010010: match <= 1'b1;
      15'b110110000010111: match <= 1'b1;
      15'b110110010111001: match <= 1'b1;
      15'b110110010111101: match <= 1'b1;
      15'b01111010100100?: match <= 1'b1;
      15'b0001110011010??: match <= 1'b1;
      15'b0101100111101??: match <= 1'b1;
      15'b1010010101011??: match <= 1'b1;
      15'b000111100001???: match <= 1'b1;
      15'b110110101011???: match <= 1'b1;
      15'b00010010000????: match <= 1'b1;
      15'b00100000000????: match <= 1'b1;
      15'b00100001011????: match <= 1'b1;
      15'b11010011110????: match <= 1'b1;
      15'b11101100011????: match <= 1'b1;
      15'b0010111100?????: match <= 1'b1;
      15'b0101111101?????: match <= 1'b1;
      15'b1001011000?????: match <= 1'b1;
      15'b1001011111?????: match <= 1'b1;
      15'b1010110011?????: match <= 1'b1;
      15'b1010110100?????: match <= 1'b1;
      15'b001010010??????: match <= 1'b1;
      15'b001010011??????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110011100(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b011001100011101: match <= 1'b1;
      15'b111110001101???: match <= 1'b1;
      15'b01010011000????: match <= 1'b1;
      15'b11111010001????: match <= 1'b1;
      15'b0101001101?????: match <= 1'b1;
      15'b1101010110?????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110011101(input clk, input rst, input [14:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      15'b000001010111100: match <= 1'b1;
      15'b100010100011100: match <= 1'b1;
      15'b100010100011101: match <= 1'b1;
      15'b100010101001101: match <= 1'b1;
      15'b100010110010010: match <= 1'b1;
      15'b100010110100101: match <= 1'b1;
      15'b101111100010001: match <= 1'b1;
      15'b101111100100001: match <= 1'b1;
      15'b101111100110000: match <= 1'b1;
      15'b10100010011????: match <= 1'b1;
      15'b10100010101????: match <= 1'b1;
      15'b10100011100????: match <= 1'b1;
      15'b10111010000????: match <= 1'b1;
      15'b10111010110????: match <= 1'b1;
      15'b10111011100????: match <= 1'b1;
      15'b0110111100?????: match <= 1'b1;
      15'b1000011111?????: match <= 1'b1;
      15'b1100000101?????: match <= 1'b1;
      15'b1100010000?????: match <= 1'b1;
      15'b1100010001?????: match <= 1'b1;
      15'b00011111???????: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110011110(input clk, input rst, input [11:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      12'b010110100111: match <= 1'b1;
      12'b01011011110?: match <= 1'b1;
      12'b10001101110?: match <= 1'b1;
      12'b1101110011??: match <= 1'b1;
      12'b001011011???: match <= 1'b1;
      12'b101101000???: match <= 1'b1;
      12'b110111001???: match <= 1'b1;
      12'b110111010???: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110011111(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b01101110110: match <= 1'b1;
      11'b11001001100: match <= 1'b1;
      11'b0110111010?: match <= 1'b1;
      11'b0110111100?: match <= 1'b1;
      11'b0110111110?: match <= 1'b1;
      11'b100100101??: match <= 1'b1;
      11'b111010000??: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110100000(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1001001110100: match <= 1'b1;
      13'b1011101000001: match <= 1'b1;
      13'b101101000100?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110100001(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b1001101100000: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110100010(input clk, input rst, input [9:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      10'b0010001110: match <= 1'b1;
      10'b1000010100: match <= 1'b1;
      10'b1011111010: match <= 1'b1;
      10'b1011111110: match <= 1'b1;
      10'b100001000?: match <= 1'b1;
      10'b110001110?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110100011(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b00101000001: match <= 1'b1;
      11'b01000010110: match <= 1'b1;
      11'b0010001000?: match <= 1'b1;
      11'b0100001010?: match <= 1'b1;
      11'b0110110010?: match <= 1'b1;
      11'b1110010110?: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110101001(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0100010100110: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110101011(input clk, input rst, input [12:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      13'b0101101001001: match <= 1'b1;
      13'b1110111000???: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110110001(input clk, input rst, input [10:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      11'b00010011001: match <= 1'b1;
      11'b00100111100: match <= 1'b1;
      11'b00110000111: match <= 1'b1;
      11'b11110100001: match <= 1'b1;
      11'b01100111???: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110111001(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0011010: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110111011(input clk, input rst, input [8:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      9'b000010011: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110111110(input clk, input rst, input [5:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      6'b000000: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module table_110111111(input clk, input rst, input [6:0] addr, output reg match);
  always@(posedge clk) begin
    casex (addr)
      7'b0101001: match <= 1'b1;
      7'b0101101: match <= 1'b1;
      7'b1111110: match <= 1'b1;
      default: match <= 1'b0;
    endcase

    if(rst)
      match <= 1'b0;
  end
endmodule

module firewall(input wire clk, input wire rst, input wire [31:0] addr,
                input wire valid, output reg match, output reg done);
  reg [31:0] addr_r;
  reg        valid_r;
  reg        match_n;

  wire out_000000010;
  table_000000010 m_000000010 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_000000010));
  wire out_000000100;
  table_000000100 m_000000100 (.clk(clk), .rst(rst), .addr(addr[22:9]), .match(out_000000100));
  wire out_000001011;
  table_000001011 m_000001011 (.clk(clk), .rst(rst), .addr(addr[22:9]), .match(out_000001011));
  wire out_000110001;
  table_000110001 m_000110001 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_000110001));
  wire out_000110110;
  table_000110110 m_000110110 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_000110110));
  wire out_000110111;
  table_000110111 m_000110111 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_000110111));
  wire out_000111110;
  table_000111110 m_000111110 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_000111110));
  wire out_001001000;
  table_001001000 m_001001000 (.clk(clk), .rst(rst), .addr(addr[22:11]), .match(out_001001000));
  wire out_001001011;
  table_001001011 m_001001011 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_001001011));
  wire out_001010010;
  table_001010010 m_001010010 (.clk(clk), .rst(rst), .addr(addr[22:11]), .match(out_001010010));
  wire out_001010100;
  table_001010100 m_001010100 (.clk(clk), .rst(rst), .addr(addr[22:13]), .match(out_001010100));
  wire out_001010101;
  table_001010101 m_001010101 (.clk(clk), .rst(rst), .addr(addr[22:20]), .match(out_001010101));
  wire out_001010111;
  table_001010111 m_001010111 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_001010111));
  wire out_001011010;
  table_001011010 m_001011010 (.clk(clk), .rst(rst), .addr(addr[22:9]), .match(out_001011010));
  wire out_001011011;
  table_001011011 m_001011011 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_001011011));
  wire out_001011100;
  table_001011100 m_001011100 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_001011100));
  wire out_001011101;
  table_001011101 m_001011101 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_001011101));
  wire out_001100011;
  table_001100011 m_001100011 (.clk(clk), .rst(rst), .addr(addr[22:13]), .match(out_001100011));
  wire out_001110100;
  table_001110100 m_001110100 (.clk(clk), .rst(rst), .addr(addr[22:17]), .match(out_001110100));
  wire out_001110111;
  table_001110111 m_001110111 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_001110111));
  wire out_001111001;
  table_001111001 m_001111001 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_001111001));
  wire out_001111010;
  table_001111010 m_001111010 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_001111010));
  wire out_001111110;
  table_001111110 m_001111110 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_001111110));
  wire out_010000000;
  table_010000000 m_010000000 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_010000000));
  wire out_010000001;
  table_010000001 m_010000001 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_010000001));
  wire out_010000010;
  table_010000010 m_010000010 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_010000010));
  wire out_010000011;
  table_010000011 m_010000011 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_010000011));
  wire out_010000111;
  table_010000111 m_010000111 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_010000111));
  wire out_010001000;
  table_010001000 m_010001000 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_010001000));
  wire out_010001010;
  table_010001010 m_010001010 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_010001010));
  wire out_010010000;
  table_010010000 m_010010000 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_010010000));
  wire out_010010100;
  table_010010100 m_010010100 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_010010100));
  wire out_010011001;
  table_010011001 m_010011001 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_010011001));
  wire out_010011010;
  table_010011010 m_010011010 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_010011010));
  wire out_010100111;
  table_010100111 m_010100111 (.clk(clk), .rst(rst), .addr(addr[22:14]), .match(out_010100111));
  wire out_010101000;
  table_010101000 m_010101000 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_010101000));
  wire out_010101001;
  table_010101001 m_010101001 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_010101001));
  wire out_010101010;
  table_010101010 m_010101010 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_010101010));
  wire out_010101011;
  table_010101011 m_010101011 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_010101011));
  wire out_010101100;
  table_010101100 m_010101100 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_010101100));
  wire out_010110001;
  table_010110001 m_010110001 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_010110001));
  wire out_010110010;
  table_010110010 m_010110010 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_010110010));
  wire out_010110111;
  table_010110111 m_010110111 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_010110111));
  wire out_010111000;
  table_010111000 m_010111000 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_010111000));
  wire out_010111010;
  table_010111010 m_010111010 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_010111010));
  wire out_010111101;
  table_010111101 m_010111101 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_010111101));
  wire out_011000000;
  table_011000000 m_011000000 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_011000000));
  wire out_011001010;
  table_011001010 m_011001010 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_011001010));
  wire out_011001011;
  table_011001011 m_011001011 (.clk(clk), .rst(rst), .addr(addr[22:13]), .match(out_011001011));
  wire out_011001101;
  table_011001101 m_011001101 (.clk(clk), .rst(rst), .addr(addr[22:13]), .match(out_011001101));
  wire out_011001110;
  table_011001110 m_011001110 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_011001110));
  wire out_011001111;
  table_011001111 m_011001111 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_011001111));
  wire out_011010001;
  table_011010001 m_011010001 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_011010001));
  wire out_011010100;
  table_011010100 m_011010100 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_011010100));
  wire out_011010111;
  table_011010111 m_011010111 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_011010111));
  wire out_011011100;
  table_011011100 m_011011100 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_011011100));
  wire out_011011111;
  table_011011111 m_011011111 (.clk(clk), .rst(rst), .addr(addr[22:13]), .match(out_011011111));
  wire out_011100011;
  table_011100011 m_011100011 (.clk(clk), .rst(rst), .addr(addr[22:13]), .match(out_011100011));
  wire out_011101001;
  table_011101001 m_011101001 (.clk(clk), .rst(rst), .addr(addr[22:17]), .match(out_011101001));
  wire out_011101010;
  table_011101010 m_011101010 (.clk(clk), .rst(rst), .addr(addr[22:15]), .match(out_011101010));
  wire out_011101110;
  table_011101110 m_011101110 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_011101110));
  wire out_011101111;
  table_011101111 m_011101111 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_011101111));
  wire out_011110000;
  table_011110000 m_011110000 (.clk(clk), .rst(rst), .addr(addr[22:17]), .match(out_011110000));
  wire out_011110100;
  table_011110100 m_011110100 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_011110100));
  wire out_011110101;
  table_011110101 m_011110101 (.clk(clk), .rst(rst), .addr(addr[22:14]), .match(out_011110101));
  wire out_011110111;
  table_011110111 m_011110111 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_011110111));
  wire out_011111000;
  table_011111000 m_011111000 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_011111000));
  wire out_011111001;
  table_011111001 m_011111001 (.clk(clk), .rst(rst), .addr(addr[22:14]), .match(out_011111001));
  wire out_011111010;
  table_011111010 m_011111010 (.clk(clk), .rst(rst), .addr(addr[22:14]), .match(out_011111010));
  wire out_011111011;
  table_011111011 m_011111011 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_011111011));
  wire out_100000000;
  table_100000000 m_100000000 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100000000));
  wire out_100000100;
  table_100000100 m_100000100 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100000100));
  wire out_100000101;
  table_100000101 m_100000101 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100000101));
  wire out_100000110;
  table_100000110 m_100000110 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_100000110));
  wire out_100000111;
  table_100000111 m_100000111 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100000111));
  wire out_100001001;
  table_100001001 m_100001001 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_100001001));
  wire out_100001100;
  table_100001100 m_100001100 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100001100));
  wire out_100001101;
  table_100001101 m_100001101 (.clk(clk), .rst(rst), .addr(addr[22:14]), .match(out_100001101));
  wire out_100010010;
  table_100010010 m_100010010 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100010010));
  wire out_100010011;
  table_100010011 m_100010011 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100010011));
  wire out_100010100;
  table_100010100 m_100010100 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_100010100));
  wire out_100010101;
  table_100010101 m_100010101 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_100010101));
  wire out_100010110;
  table_100010110 m_100010110 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100010110));
  wire out_100010111;
  table_100010111 m_100010111 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100010111));
  wire out_100011000;
  table_100011000 m_100011000 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_100011000));
  wire out_100011001;
  table_100011001 m_100011001 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100011001));
  wire out_100011010;
  table_100011010 m_100011010 (.clk(clk), .rst(rst), .addr(addr[22:9]), .match(out_100011010));
  wire out_100011011;
  table_100011011 m_100011011 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_100011011));
  wire out_100011100;
  table_100011100 m_100011100 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100011100));
  wire out_100011110;
  table_100011110 m_100011110 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_100011110));
  wire out_100011111;
  table_100011111 m_100011111 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100011111));
  wire out_100100011;
  table_100100011 m_100100011 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100100011));
  wire out_100100100;
  table_100100100 m_100100100 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100100100));
  wire out_100100101;
  table_100100101 m_100100101 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100100101));
  wire out_100100110;
  table_100100110 m_100100110 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_100100110));
  wire out_100101001;
  table_100101001 m_100101001 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100101001));
  wire out_100101010;
  table_100101010 m_100101010 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100101010));
  wire out_100101011;
  table_100101011 m_100101011 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100101011));
  wire out_100101100;
  table_100101100 m_100101100 (.clk(clk), .rst(rst), .addr(addr[22:15]), .match(out_100101100));
  wire out_100101101;
  table_100101101 m_100101101 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_100101101));
  wire out_100101111;
  table_100101111 m_100101111 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100101111));
  wire out_100110000;
  table_100110000 m_100110000 (.clk(clk), .rst(rst), .addr(addr[22:9]), .match(out_100110000));
  wire out_100110001;
  table_100110001 m_100110001 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100110001));
  wire out_100110010;
  table_100110010 m_100110010 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100110010));
  wire out_100110110;
  table_100110110 m_100110110 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100110110));
  wire out_100110111;
  table_100110111 m_100110111 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100110111));
  wire out_100111000;
  table_100111000 m_100111000 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100111000));
  wire out_100111001;
  table_100111001 m_100111001 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_100111001));
  wire out_100111010;
  table_100111010 m_100111010 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100111010));
  wire out_100111011;
  table_100111011 m_100111011 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100111011));
  wire out_100111100;
  table_100111100 m_100111100 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100111100));
  wire out_100111101;
  table_100111101 m_100111101 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100111101));
  wire out_100111110;
  table_100111110 m_100111110 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100111110));
  wire out_100111111;
  table_100111111 m_100111111 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_100111111));
  wire out_101000000;
  table_101000000 m_101000000 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_101000000));
  wire out_101000001;
  table_101000001 m_101000001 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_101000001));
  wire out_101000010;
  table_101000010 m_101000010 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_101000010));
  wire out_101000101;
  table_101000101 m_101000101 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_101000101));
  wire out_101000110;
  table_101000110 m_101000110 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_101000110));
  wire out_101000111;
  table_101000111 m_101000111 (.clk(clk), .rst(rst), .addr(addr[22:13]), .match(out_101000111));
  wire out_101001000;
  table_101001000 m_101001000 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_101001000));
  wire out_101001001;
  table_101001001 m_101001001 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_101001001));
  wire out_101001010;
  table_101001010 m_101001010 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_101001010));
  wire out_101001011;
  table_101001011 m_101001011 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_101001011));
  wire out_101001100;
  table_101001100 m_101001100 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_101001100));
  wire out_101001110;
  table_101001110 m_101001110 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_101001110));
  wire out_101001111;
  table_101001111 m_101001111 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_101001111));
  wire out_101010000;
  table_101010000 m_101010000 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_101010000));
  wire out_101010001;
  table_101010001 m_101010001 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_101010001));
  wire out_101010011;
  table_101010011 m_101010011 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_101010011));
  wire out_101010100;
  table_101010100 m_101010100 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_101010100));
  wire out_101010101;
  table_101010101 m_101010101 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_101010101));
  wire out_101010110;
  table_101010110 m_101010110 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_101010110));
  wire out_101011110;
  table_101011110 m_101011110 (.clk(clk), .rst(rst), .addr(addr[22:14]), .match(out_101011110));
  wire out_101100000;
  table_101100000 m_101100000 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_101100000));
  wire out_101100001;
  table_101100001 m_101100001 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_101100001));
  wire out_101100011;
  table_101100011 m_101100011 (.clk(clk), .rst(rst), .addr(addr[22:11]), .match(out_101100011));
  wire out_101100101;
  table_101100101 m_101100101 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_101100101));
  wire out_101100110;
  table_101100110 m_101100110 (.clk(clk), .rst(rst), .addr(addr[22:15]), .match(out_101100110));
  wire out_101101001;
  table_101101001 m_101101001 (.clk(clk), .rst(rst), .addr(addr[22:14]), .match(out_101101001));
  wire out_101101011;
  table_101101011 m_101101011 (.clk(clk), .rst(rst), .addr(addr[22:11]), .match(out_101101011));
  wire out_101110010;
  table_101110010 m_101110010 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_101110010));
  wire out_101110011;
  table_101110011 m_101110011 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_101110011));
  wire out_101110100;
  table_101110100 m_101110100 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_101110100));
  wire out_101110101;
  table_101110101 m_101110101 (.clk(clk), .rst(rst), .addr(addr[22:14]), .match(out_101110101));
  wire out_101111001;
  table_101111001 m_101111001 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_101111001));
  wire out_101111100;
  table_101111100 m_101111100 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_101111100));
  wire out_101111101;
  table_101111101 m_101111101 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_101111101));
  wire out_110000000;
  table_110000000 m_110000000 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110000000));
  wire out_110000001;
  table_110000001 m_110000001 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110000001));
  wire out_110000010;
  table_110000010 m_110000010 (.clk(clk), .rst(rst), .addr(addr[22:9]), .match(out_110000010));
  wire out_110000011;
  table_110000011 m_110000011 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110000011));
  wire out_110000100;
  table_110000100 m_110000100 (.clk(clk), .rst(rst), .addr(addr[22:9]), .match(out_110000100));
  wire out_110000101;
  table_110000101 m_110000101 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110000101));
  wire out_110000111;
  table_110000111 m_110000111 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110000111));
  wire out_110001000;
  table_110001000 m_110001000 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110001000));
  wire out_110001001;
  table_110001001 m_110001001 (.clk(clk), .rst(rst), .addr(addr[22:14]), .match(out_110001001));
  wire out_110001011;
  table_110001011 m_110001011 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_110001011));
  wire out_110001100;
  table_110001100 m_110001100 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110001100));
  wire out_110001101;
  table_110001101 m_110001101 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110001101));
  wire out_110001110;
  table_110001110 m_110001110 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110001110));
  wire out_110001111;
  table_110001111 m_110001111 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110001111));
  wire out_110010000;
  table_110010000 m_110010000 (.clk(clk), .rst(rst), .addr(addr[22:9]), .match(out_110010000));
  wire out_110010001;
  table_110010001 m_110010001 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_110010001));
  wire out_110010011;
  table_110010011 m_110010011 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_110010011));
  wire out_110010100;
  table_110010100 m_110010100 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110010100));
  wire out_110010101;
  table_110010101 m_110010101 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_110010101));
  wire out_110010110;
  table_110010110 m_110010110 (.clk(clk), .rst(rst), .addr(addr[22:9]), .match(out_110010110));
  wire out_110010111;
  table_110010111 m_110010111 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_110010111));
  wire out_110011000;
  table_110011000 m_110011000 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110011000));
  wire out_110011001;
  table_110011001 m_110011001 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110011001));
  wire out_110011011;
  table_110011011 m_110011011 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110011011));
  wire out_110011100;
  table_110011100 m_110011100 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110011100));
  wire out_110011101;
  table_110011101 m_110011101 (.clk(clk), .rst(rst), .addr(addr[22:8]), .match(out_110011101));
  wire out_110011110;
  table_110011110 m_110011110 (.clk(clk), .rst(rst), .addr(addr[22:11]), .match(out_110011110));
  wire out_110011111;
  table_110011111 m_110011111 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_110011111));
  wire out_110100000;
  table_110100000 m_110100000 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_110100000));
  wire out_110100001;
  table_110100001 m_110100001 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_110100001));
  wire out_110100010;
  table_110100010 m_110100010 (.clk(clk), .rst(rst), .addr(addr[22:13]), .match(out_110100010));
  wire out_110100011;
  table_110100011 m_110100011 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_110100011));
  wire out_110101001;
  table_110101001 m_110101001 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_110101001));
  wire out_110101011;
  table_110101011 m_110101011 (.clk(clk), .rst(rst), .addr(addr[22:10]), .match(out_110101011));
  wire out_110110001;
  table_110110001 m_110110001 (.clk(clk), .rst(rst), .addr(addr[22:12]), .match(out_110110001));
  wire out_110111001;
  table_110111001 m_110111001 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_110111001));
  wire out_110111011;
  table_110111011 m_110111011 (.clk(clk), .rst(rst), .addr(addr[22:14]), .match(out_110111011));
  wire out_110111110;
  table_110111110 m_110111110 (.clk(clk), .rst(rst), .addr(addr[22:17]), .match(out_110111110));
  wire out_110111111;
  table_110111111 m_110111111 (.clk(clk), .rst(rst), .addr(addr[22:16]), .match(out_110111111));

  always@(*)
    case (addr_r[31:23])
      9'b000000010: match_n = out_000000010;
      9'b000000100: match_n = out_000000100;
      9'b000001011: match_n = out_000001011;
      9'b000110001: match_n = out_000110001;
      9'b000110110: match_n = out_000110110;
      9'b000110111: match_n = out_000110111;
      9'b000111110: match_n = out_000111110;
      9'b001001000: match_n = out_001001000;
      9'b001001011: match_n = out_001001011;
      9'b001010010: match_n = out_001010010;
      9'b001010100: match_n = out_001010100;
      9'b001010101: match_n = out_001010101;
      9'b001010111: match_n = out_001010111;
      9'b001011010: match_n = out_001011010;
      9'b001011011: match_n = out_001011011;
      9'b001011100: match_n = out_001011100;
      9'b001011101: match_n = out_001011101;
      9'b001100011: match_n = out_001100011;
      9'b001110100: match_n = out_001110100;
      9'b001110111: match_n = out_001110111;
      9'b001111001: match_n = out_001111001;
      9'b001111010: match_n = out_001111010;
      9'b001111110: match_n = out_001111110;
      9'b010000000: match_n = out_010000000;
      9'b010000001: match_n = out_010000001;
      9'b010000010: match_n = out_010000010;
      9'b010000011: match_n = out_010000011;
      9'b010000111: match_n = out_010000111;
      9'b010001000: match_n = out_010001000;
      9'b010001010: match_n = out_010001010;
      9'b010010000: match_n = out_010010000;
      9'b010010100: match_n = out_010010100;
      9'b010011001: match_n = out_010011001;
      9'b010011010: match_n = out_010011010;
      9'b010100111: match_n = out_010100111;
      9'b010101000: match_n = out_010101000;
      9'b010101001: match_n = out_010101001;
      9'b010101010: match_n = out_010101010;
      9'b010101011: match_n = out_010101011;
      9'b010101100: match_n = out_010101100;
      9'b010110001: match_n = out_010110001;
      9'b010110010: match_n = out_010110010;
      9'b010110111: match_n = out_010110111;
      9'b010111000: match_n = out_010111000;
      9'b010111010: match_n = out_010111010;
      9'b010111101: match_n = out_010111101;
      9'b011000000: match_n = out_011000000;
      9'b011001010: match_n = out_011001010;
      9'b011001011: match_n = out_011001011;
      9'b011001101: match_n = out_011001101;
      9'b011001110: match_n = out_011001110;
      9'b011001111: match_n = out_011001111;
      9'b011010001: match_n = out_011010001;
      9'b011010100: match_n = out_011010100;
      9'b011010111: match_n = out_011010111;
      9'b011011100: match_n = out_011011100;
      9'b011011111: match_n = out_011011111;
      9'b011100011: match_n = out_011100011;
      9'b011101001: match_n = out_011101001;
      9'b011101010: match_n = out_011101010;
      9'b011101110: match_n = out_011101110;
      9'b011101111: match_n = out_011101111;
      9'b011110000: match_n = out_011110000;
      9'b011110100: match_n = out_011110100;
      9'b011110101: match_n = out_011110101;
      9'b011110111: match_n = out_011110111;
      9'b011111000: match_n = out_011111000;
      9'b011111001: match_n = out_011111001;
      9'b011111010: match_n = out_011111010;
      9'b011111011: match_n = out_011111011;
      9'b100000000: match_n = out_100000000;
      9'b100000100: match_n = out_100000100;
      9'b100000101: match_n = out_100000101;
      9'b100000110: match_n = out_100000110;
      9'b100000111: match_n = out_100000111;
      9'b100001001: match_n = out_100001001;
      9'b100001100: match_n = out_100001100;
      9'b100001101: match_n = out_100001101;
      9'b100010010: match_n = out_100010010;
      9'b100010011: match_n = out_100010011;
      9'b100010100: match_n = out_100010100;
      9'b100010101: match_n = out_100010101;
      9'b100010110: match_n = out_100010110;
      9'b100010111: match_n = out_100010111;
      9'b100011000: match_n = out_100011000;
      9'b100011001: match_n = out_100011001;
      9'b100011010: match_n = out_100011010;
      9'b100011011: match_n = out_100011011;
      9'b100011100: match_n = out_100011100;
      9'b100011110: match_n = out_100011110;
      9'b100011111: match_n = out_100011111;
      9'b100100011: match_n = out_100100011;
      9'b100100100: match_n = out_100100100;
      9'b100100101: match_n = out_100100101;
      9'b100100110: match_n = out_100100110;
      9'b100101001: match_n = out_100101001;
      9'b100101010: match_n = out_100101010;
      9'b100101011: match_n = out_100101011;
      9'b100101100: match_n = out_100101100;
      9'b100101101: match_n = out_100101101;
      9'b100101111: match_n = out_100101111;
      9'b100110000: match_n = out_100110000;
      9'b100110001: match_n = out_100110001;
      9'b100110010: match_n = out_100110010;
      9'b100110110: match_n = out_100110110;
      9'b100110111: match_n = out_100110111;
      9'b100111000: match_n = out_100111000;
      9'b100111001: match_n = out_100111001;
      9'b100111010: match_n = out_100111010;
      9'b100111011: match_n = out_100111011;
      9'b100111100: match_n = out_100111100;
      9'b100111101: match_n = out_100111101;
      9'b100111110: match_n = out_100111110;
      9'b100111111: match_n = out_100111111;
      9'b101000000: match_n = out_101000000;
      9'b101000001: match_n = out_101000001;
      9'b101000010: match_n = out_101000010;
      9'b101000101: match_n = out_101000101;
      9'b101000110: match_n = out_101000110;
      9'b101000111: match_n = out_101000111;
      9'b101001000: match_n = out_101001000;
      9'b101001001: match_n = out_101001001;
      9'b101001010: match_n = out_101001010;
      9'b101001011: match_n = out_101001011;
      9'b101001100: match_n = out_101001100;
      9'b101001110: match_n = out_101001110;
      9'b101001111: match_n = out_101001111;
      9'b101010000: match_n = out_101010000;
      9'b101010001: match_n = out_101010001;
      9'b101010011: match_n = out_101010011;
      9'b101010100: match_n = out_101010100;
      9'b101010101: match_n = out_101010101;
      9'b101010110: match_n = out_101010110;
      9'b101011110: match_n = out_101011110;
      9'b101100000: match_n = out_101100000;
      9'b101100001: match_n = out_101100001;
      9'b101100011: match_n = out_101100011;
      9'b101100101: match_n = out_101100101;
      9'b101100110: match_n = out_101100110;
      9'b101101001: match_n = out_101101001;
      9'b101101011: match_n = out_101101011;
      9'b101110010: match_n = out_101110010;
      9'b101110011: match_n = out_101110011;
      9'b101110100: match_n = out_101110100;
      9'b101110101: match_n = out_101110101;
      9'b101111001: match_n = out_101111001;
      9'b101111100: match_n = out_101111100;
      9'b101111101: match_n = out_101111101;
      9'b110000000: match_n = out_110000000;
      9'b110000001: match_n = out_110000001;
      9'b110000010: match_n = out_110000010;
      9'b110000011: match_n = out_110000011;
      9'b110000100: match_n = out_110000100;
      9'b110000101: match_n = out_110000101;
      9'b110000111: match_n = out_110000111;
      9'b110001000: match_n = out_110001000;
      9'b110001001: match_n = out_110001001;
      9'b110001011: match_n = out_110001011;
      9'b110001100: match_n = out_110001100;
      9'b110001101: match_n = out_110001101;
      9'b110001110: match_n = out_110001110;
      9'b110001111: match_n = out_110001111;
      9'b110010000: match_n = out_110010000;
      9'b110010001: match_n = out_110010001;
      9'b110010011: match_n = out_110010011;
      9'b110010100: match_n = out_110010100;
      9'b110010101: match_n = out_110010101;
      9'b110010110: match_n = out_110010110;
      9'b110010111: match_n = out_110010111;
      9'b110011000: match_n = out_110011000;
      9'b110011001: match_n = out_110011001;
      9'b110011011: match_n = out_110011011;
      9'b110011100: match_n = out_110011100;
      9'b110011101: match_n = out_110011101;
      9'b110011110: match_n = out_110011110;
      9'b110011111: match_n = out_110011111;
      9'b110100000: match_n = out_110100000;
      9'b110100001: match_n = out_110100001;
      9'b110100010: match_n = out_110100010;
      9'b110100011: match_n = out_110100011;
      9'b110101001: match_n = out_110101001;
      9'b110101011: match_n = out_110101011;
      9'b110110001: match_n = out_110110001;
      9'b110111001: match_n = out_110111001;
      9'b110111011: match_n = out_110111011;
      9'b110111110: match_n = out_110111110;
      9'b110111111: match_n = out_110111111;
      default: match_n = 1'b0;
    endcase

  always@(posedge clk) begin
    addr_r  <= addr;
    valid_r <= valid;
    match   <= (match || match_n) && !valid;
    done    <= (done  || valid_r) && !valid;

    if(rst) begin
      match   <= 1'b0;
      done    <= 1'b0;
      valid_r <= 1'b0;
    end
  end
endmodule

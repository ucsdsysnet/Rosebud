`include "struct_s.sv"
module string_matcher (
    clk,
    rst,
    in_data,
    in_valid,
    init,
    in_last,
    in_strb,
    in_ready,
    out_data,
    out_valid,
    out_almost_full,
    out_last
);

input clk;
input rst;
input [255:0] in_data;
input in_valid;
input init;
input in_last;
input [7:0] in_strb;
output logic in_ready;
output logic [127:0] out_data;
output logic out_valid;
output logic out_last;
input out_almost_full;

logic [255:0] in_data_r1;
logic [255:0] in_data_r2;
logic         in_valid_r1;
logic         in_valid_r2;
logic         init_r1;
logic         init_r2;
logic         in_last_r1;
logic         in_last_r2;
logic [7:0]   in_strb_r1;
logic [7:0]   in_strb_r2;

logic [RID_WIDTH-1:0] hash_out_0_0;
logic hash_out_valid_filter_0_0;
rule_s_t din_0_0;
rule_s_t din_0_0_r1;
rule_s_t din_0_0_r2;
logic din_valid_0_0;
logic din_valid_0_0_r1;
logic din_valid_0_0_r2;
logic din_almost_full_0_0;
logic [RID_WIDTH-1:0] hash_out_0_1;
logic hash_out_valid_filter_0_1;
rule_s_t din_0_1;
rule_s_t din_0_1_r1;
rule_s_t din_0_1_r2;
logic din_valid_0_1;
logic din_valid_0_1_r1;
logic din_valid_0_1_r2;
logic din_almost_full_0_1;
logic [RID_WIDTH-1:0] hash_out_0_2;
logic hash_out_valid_filter_0_2;
rule_s_t din_0_2;
rule_s_t din_0_2_r1;
rule_s_t din_0_2_r2;
logic din_valid_0_2;
logic din_valid_0_2_r1;
logic din_valid_0_2_r2;
logic din_almost_full_0_2;
logic [RID_WIDTH-1:0] hash_out_0_3;
logic hash_out_valid_filter_0_3;
rule_s_t din_0_3;
rule_s_t din_0_3_r1;
rule_s_t din_0_3_r2;
logic din_valid_0_3;
logic din_valid_0_3_r1;
logic din_valid_0_3_r2;
logic din_almost_full_0_3;
logic [RID_WIDTH-1:0] hash_out_0_4;
logic hash_out_valid_filter_0_4;
rule_s_t din_0_4;
rule_s_t din_0_4_r1;
rule_s_t din_0_4_r2;
logic din_valid_0_4;
logic din_valid_0_4_r1;
logic din_valid_0_4_r2;
logic din_almost_full_0_4;
logic [RID_WIDTH-1:0] hash_out_0_5;
logic hash_out_valid_filter_0_5;
rule_s_t din_0_5;
rule_s_t din_0_5_r1;
rule_s_t din_0_5_r2;
logic din_valid_0_5;
logic din_valid_0_5_r1;
logic din_valid_0_5_r2;
logic din_almost_full_0_5;
logic [RID_WIDTH-1:0] hash_out_0_6;
logic hash_out_valid_filter_0_6;
rule_s_t din_0_6;
rule_s_t din_0_6_r1;
rule_s_t din_0_6_r2;
logic din_valid_0_6;
logic din_valid_0_6_r1;
logic din_valid_0_6_r2;
logic din_almost_full_0_6;
logic [RID_WIDTH-1:0] hash_out_0_7;
logic hash_out_valid_filter_0_7;
rule_s_t din_0_7;
rule_s_t din_0_7_r1;
rule_s_t din_0_7_r2;
logic din_valid_0_7;
logic din_valid_0_7_r1;
logic din_valid_0_7_r2;
logic din_almost_full_0_7;

rule_s_t din_0_8_r2;
logic din_valid_0_8_r2 = 1'b0;
logic din_almost_full_0_8;
assign din_0_8_r2.data   = 0;
assign din_0_8_r2.last   = 1'b0;
assign din_0_8_r2.bucket = 0;
rule_s_t din_0_9_r2;
logic din_valid_0_9_r2 = 1'b0;
logic din_almost_full_0_9;
assign din_0_9_r2.data   = 0;
assign din_0_9_r2.last   = 1'b0;
assign din_0_9_r2.bucket = 0;
rule_s_t din_0_10_r2;
logic din_valid_0_10_r2 = 1'b0;
logic din_almost_full_0_10;
assign din_0_10_r2.data   = 0;
assign din_0_10_r2.last   = 1'b0;
assign din_0_10_r2.bucket = 0;
rule_s_t din_0_11_r2;
logic din_valid_0_11_r2 = 1'b0;
logic din_almost_full_0_11;
assign din_0_11_r2.data   = 0;
assign din_0_11_r2.last   = 1'b0;
assign din_0_11_r2.bucket = 0;
rule_s_t din_0_12_r2;
logic din_valid_0_12_r2 = 1'b0;
logic din_almost_full_0_12;
assign din_0_12_r2.data   = 0;
assign din_0_12_r2.last   = 1'b0;
assign din_0_12_r2.bucket = 0;
rule_s_t din_0_13_r2;
logic din_valid_0_13_r2 = 1'b0;
logic din_almost_full_0_13;
assign din_0_13_r2.data   = 0;
assign din_0_13_r2.last   = 1'b0;
assign din_0_13_r2.bucket = 0;
rule_s_t din_0_14_r2;
logic din_valid_0_14_r2 = 1'b0;
logic din_almost_full_0_14;
assign din_0_14_r2.data   = 0;
assign din_0_14_r2.last   = 1'b0;
assign din_0_14_r2.bucket = 0;
rule_s_t din_0_15_r2;
logic din_valid_0_15_r2 = 1'b0;
logic din_almost_full_0_15;
assign din_0_15_r2.data   = 0;
assign din_0_15_r2.last   = 1'b0;
assign din_0_15_r2.bucket = 0;
rule_s_t din_0_16_r2;
logic din_valid_0_16_r2 = 1'b0;
logic din_almost_full_0_16;
assign din_0_16_r2.data   = 0;
assign din_0_16_r2.last   = 1'b0;
assign din_0_16_r2.bucket = 0;
rule_s_t din_0_17_r2;
logic din_valid_0_17_r2 = 1'b0;
logic din_almost_full_0_17;
assign din_0_17_r2.data   = 0;
assign din_0_17_r2.last   = 1'b0;
assign din_0_17_r2.bucket = 0;
rule_s_t din_0_18_r2;
logic din_valid_0_18_r2 = 1'b0;
logic din_almost_full_0_18;
assign din_0_18_r2.data   = 0;
assign din_0_18_r2.last   = 1'b0;
assign din_0_18_r2.bucket = 0;
rule_s_t din_0_19_r2;
logic din_valid_0_19_r2 = 1'b0;
logic din_almost_full_0_19;
assign din_0_19_r2.data   = 0;
assign din_0_19_r2.last   = 1'b0;
assign din_0_19_r2.bucket = 0;
rule_s_t din_0_20_r2;
logic din_valid_0_20_r2 = 1'b0;
logic din_almost_full_0_20;
assign din_0_20_r2.data   = 0;
assign din_0_20_r2.last   = 1'b0;
assign din_0_20_r2.bucket = 0;
rule_s_t din_0_21_r2;
logic din_valid_0_21_r2 = 1'b0;
logic din_almost_full_0_21;
assign din_0_21_r2.data   = 0;
assign din_0_21_r2.last   = 1'b0;
assign din_0_21_r2.bucket = 0;
rule_s_t din_0_22_r2;
logic din_valid_0_22_r2 = 1'b0;
logic din_almost_full_0_22;
assign din_0_22_r2.data   = 0;
assign din_0_22_r2.last   = 1'b0;
assign din_0_22_r2.bucket = 0;
rule_s_t din_0_23_r2;
logic din_valid_0_23_r2 = 1'b0;
logic din_almost_full_0_23;
assign din_0_23_r2.data   = 0;
assign din_0_23_r2.last   = 1'b0;
assign din_0_23_r2.bucket = 0;
rule_s_t din_0_24_r2;
logic din_valid_0_24_r2 = 1'b0;
logic din_almost_full_0_24;
assign din_0_24_r2.data   = 0;
assign din_0_24_r2.last   = 1'b0;
assign din_0_24_r2.bucket = 0;
rule_s_t din_0_25_r2;
logic din_valid_0_25_r2 = 1'b0;
logic din_almost_full_0_25;
assign din_0_25_r2.data   = 0;
assign din_0_25_r2.last   = 1'b0;
assign din_0_25_r2.bucket = 0;
rule_s_t din_0_26_r2;
logic din_valid_0_26_r2 = 1'b0;
logic din_almost_full_0_26;
assign din_0_26_r2.data   = 0;
assign din_0_26_r2.last   = 1'b0;
assign din_0_26_r2.bucket = 0;
rule_s_t din_0_27_r2;
logic din_valid_0_27_r2 = 1'b0;
logic din_almost_full_0_27;
assign din_0_27_r2.data   = 0;
assign din_0_27_r2.last   = 1'b0;
assign din_0_27_r2.bucket = 0;
rule_s_t din_0_28_r2;
logic din_valid_0_28_r2 = 1'b0;
logic din_almost_full_0_28;
assign din_0_28_r2.data   = 0;
assign din_0_28_r2.last   = 1'b0;
assign din_0_28_r2.bucket = 0;
rule_s_t din_0_29_r2;
logic din_valid_0_29_r2 = 1'b0;
logic din_almost_full_0_29;
assign din_0_29_r2.data   = 0;
assign din_0_29_r2.last   = 1'b0;
assign din_0_29_r2.bucket = 0;
rule_s_t din_0_30_r2;
logic din_valid_0_30_r2 = 1'b0;
logic din_almost_full_0_30;
assign din_0_30_r2.data   = 0;
assign din_0_30_r2.last   = 1'b0;
assign din_0_30_r2.bucket = 0;
rule_s_t din_0_31_r2;
logic din_valid_0_31_r2 = 1'b0;
logic din_almost_full_0_31;
assign din_0_31_r2.data   = 0;
assign din_0_31_r2.last   = 1'b0;
assign din_0_31_r2.bucket = 0;

logic [RID_WIDTH-1:0] hash_out_1_0;
logic hash_out_valid_filter_1_0;
rule_s_t din_1_0;
rule_s_t din_1_0_r1;
rule_s_t din_1_0_r2;
logic din_valid_1_0;
logic din_valid_1_0_r1;
logic din_valid_1_0_r2;
logic din_almost_full_1_0;
logic [RID_WIDTH-1:0] hash_out_1_1;
logic hash_out_valid_filter_1_1;
rule_s_t din_1_1;
rule_s_t din_1_1_r1;
rule_s_t din_1_1_r2;
logic din_valid_1_1;
logic din_valid_1_1_r1;
logic din_valid_1_1_r2;
logic din_almost_full_1_1;
logic [RID_WIDTH-1:0] hash_out_1_2;
logic hash_out_valid_filter_1_2;
rule_s_t din_1_2;
rule_s_t din_1_2_r1;
rule_s_t din_1_2_r2;
logic din_valid_1_2;
logic din_valid_1_2_r1;
logic din_valid_1_2_r2;
logic din_almost_full_1_2;
logic [RID_WIDTH-1:0] hash_out_1_3;
logic hash_out_valid_filter_1_3;
rule_s_t din_1_3;
rule_s_t din_1_3_r1;
rule_s_t din_1_3_r2;
logic din_valid_1_3;
logic din_valid_1_3_r1;
logic din_valid_1_3_r2;
logic din_almost_full_1_3;
logic [RID_WIDTH-1:0] hash_out_1_4;
logic hash_out_valid_filter_1_4;
rule_s_t din_1_4;
rule_s_t din_1_4_r1;
rule_s_t din_1_4_r2;
logic din_valid_1_4;
logic din_valid_1_4_r1;
logic din_valid_1_4_r2;
logic din_almost_full_1_4;
logic [RID_WIDTH-1:0] hash_out_1_5;
logic hash_out_valid_filter_1_5;
rule_s_t din_1_5;
rule_s_t din_1_5_r1;
rule_s_t din_1_5_r2;
logic din_valid_1_5;
logic din_valid_1_5_r1;
logic din_valid_1_5_r2;
logic din_almost_full_1_5;
logic [RID_WIDTH-1:0] hash_out_1_6;
logic hash_out_valid_filter_1_6;
rule_s_t din_1_6;
rule_s_t din_1_6_r1;
rule_s_t din_1_6_r2;
logic din_valid_1_6;
logic din_valid_1_6_r1;
logic din_valid_1_6_r2;
logic din_almost_full_1_6;
logic [RID_WIDTH-1:0] hash_out_1_7;
logic hash_out_valid_filter_1_7;
rule_s_t din_1_7;
rule_s_t din_1_7_r1;
rule_s_t din_1_7_r2;
logic din_valid_1_7;
logic din_valid_1_7_r1;
logic din_valid_1_7_r2;
logic din_almost_full_1_7;

rule_s_t din_1_8_r2;
logic din_valid_1_8_r2 = 1'b0;
logic din_almost_full_1_8;
assign din_1_8_r2.data   = 0;
assign din_1_8_r2.last   = 1'b0;
assign din_1_8_r2.bucket = 1;
rule_s_t din_1_9_r2;
logic din_valid_1_9_r2 = 1'b0;
logic din_almost_full_1_9;
assign din_1_9_r2.data   = 0;
assign din_1_9_r2.last   = 1'b0;
assign din_1_9_r2.bucket = 1;
rule_s_t din_1_10_r2;
logic din_valid_1_10_r2 = 1'b0;
logic din_almost_full_1_10;
assign din_1_10_r2.data   = 0;
assign din_1_10_r2.last   = 1'b0;
assign din_1_10_r2.bucket = 1;
rule_s_t din_1_11_r2;
logic din_valid_1_11_r2 = 1'b0;
logic din_almost_full_1_11;
assign din_1_11_r2.data   = 0;
assign din_1_11_r2.last   = 1'b0;
assign din_1_11_r2.bucket = 1;
rule_s_t din_1_12_r2;
logic din_valid_1_12_r2 = 1'b0;
logic din_almost_full_1_12;
assign din_1_12_r2.data   = 0;
assign din_1_12_r2.last   = 1'b0;
assign din_1_12_r2.bucket = 1;
rule_s_t din_1_13_r2;
logic din_valid_1_13_r2 = 1'b0;
logic din_almost_full_1_13;
assign din_1_13_r2.data   = 0;
assign din_1_13_r2.last   = 1'b0;
assign din_1_13_r2.bucket = 1;
rule_s_t din_1_14_r2;
logic din_valid_1_14_r2 = 1'b0;
logic din_almost_full_1_14;
assign din_1_14_r2.data   = 0;
assign din_1_14_r2.last   = 1'b0;
assign din_1_14_r2.bucket = 1;
rule_s_t din_1_15_r2;
logic din_valid_1_15_r2 = 1'b0;
logic din_almost_full_1_15;
assign din_1_15_r2.data   = 0;
assign din_1_15_r2.last   = 1'b0;
assign din_1_15_r2.bucket = 1;
rule_s_t din_1_16_r2;
logic din_valid_1_16_r2 = 1'b0;
logic din_almost_full_1_16;
assign din_1_16_r2.data   = 0;
assign din_1_16_r2.last   = 1'b0;
assign din_1_16_r2.bucket = 1;
rule_s_t din_1_17_r2;
logic din_valid_1_17_r2 = 1'b0;
logic din_almost_full_1_17;
assign din_1_17_r2.data   = 0;
assign din_1_17_r2.last   = 1'b0;
assign din_1_17_r2.bucket = 1;
rule_s_t din_1_18_r2;
logic din_valid_1_18_r2 = 1'b0;
logic din_almost_full_1_18;
assign din_1_18_r2.data   = 0;
assign din_1_18_r2.last   = 1'b0;
assign din_1_18_r2.bucket = 1;
rule_s_t din_1_19_r2;
logic din_valid_1_19_r2 = 1'b0;
logic din_almost_full_1_19;
assign din_1_19_r2.data   = 0;
assign din_1_19_r2.last   = 1'b0;
assign din_1_19_r2.bucket = 1;
rule_s_t din_1_20_r2;
logic din_valid_1_20_r2 = 1'b0;
logic din_almost_full_1_20;
assign din_1_20_r2.data   = 0;
assign din_1_20_r2.last   = 1'b0;
assign din_1_20_r2.bucket = 1;
rule_s_t din_1_21_r2;
logic din_valid_1_21_r2 = 1'b0;
logic din_almost_full_1_21;
assign din_1_21_r2.data   = 0;
assign din_1_21_r2.last   = 1'b0;
assign din_1_21_r2.bucket = 1;
rule_s_t din_1_22_r2;
logic din_valid_1_22_r2 = 1'b0;
logic din_almost_full_1_22;
assign din_1_22_r2.data   = 0;
assign din_1_22_r2.last   = 1'b0;
assign din_1_22_r2.bucket = 1;
rule_s_t din_1_23_r2;
logic din_valid_1_23_r2 = 1'b0;
logic din_almost_full_1_23;
assign din_1_23_r2.data   = 0;
assign din_1_23_r2.last   = 1'b0;
assign din_1_23_r2.bucket = 1;
rule_s_t din_1_24_r2;
logic din_valid_1_24_r2 = 1'b0;
logic din_almost_full_1_24;
assign din_1_24_r2.data   = 0;
assign din_1_24_r2.last   = 1'b0;
assign din_1_24_r2.bucket = 1;
rule_s_t din_1_25_r2;
logic din_valid_1_25_r2 = 1'b0;
logic din_almost_full_1_25;
assign din_1_25_r2.data   = 0;
assign din_1_25_r2.last   = 1'b0;
assign din_1_25_r2.bucket = 1;
rule_s_t din_1_26_r2;
logic din_valid_1_26_r2 = 1'b0;
logic din_almost_full_1_26;
assign din_1_26_r2.data   = 0;
assign din_1_26_r2.last   = 1'b0;
assign din_1_26_r2.bucket = 1;
rule_s_t din_1_27_r2;
logic din_valid_1_27_r2 = 1'b0;
logic din_almost_full_1_27;
assign din_1_27_r2.data   = 0;
assign din_1_27_r2.last   = 1'b0;
assign din_1_27_r2.bucket = 1;
rule_s_t din_1_28_r2;
logic din_valid_1_28_r2 = 1'b0;
logic din_almost_full_1_28;
assign din_1_28_r2.data   = 0;
assign din_1_28_r2.last   = 1'b0;
assign din_1_28_r2.bucket = 1;
rule_s_t din_1_29_r2;
logic din_valid_1_29_r2 = 1'b0;
logic din_almost_full_1_29;
assign din_1_29_r2.data   = 0;
assign din_1_29_r2.last   = 1'b0;
assign din_1_29_r2.bucket = 1;
rule_s_t din_1_30_r2;
logic din_valid_1_30_r2 = 1'b0;
logic din_almost_full_1_30;
assign din_1_30_r2.data   = 0;
assign din_1_30_r2.last   = 1'b0;
assign din_1_30_r2.bucket = 1;
rule_s_t din_1_31_r2;
logic din_valid_1_31_r2 = 1'b0;
logic din_almost_full_1_31;
assign din_1_31_r2.data   = 0;
assign din_1_31_r2.last   = 1'b0;
assign din_1_31_r2.bucket = 1;

logic [RID_WIDTH-1:0] hash_out_2_0;
logic hash_out_valid_filter_2_0;
rule_s_t din_2_0;
rule_s_t din_2_0_r1;
rule_s_t din_2_0_r2;
logic din_valid_2_0;
logic din_valid_2_0_r1;
logic din_valid_2_0_r2;
logic din_almost_full_2_0;
logic [RID_WIDTH-1:0] hash_out_2_1;
logic hash_out_valid_filter_2_1;
rule_s_t din_2_1;
rule_s_t din_2_1_r1;
rule_s_t din_2_1_r2;
logic din_valid_2_1;
logic din_valid_2_1_r1;
logic din_valid_2_1_r2;
logic din_almost_full_2_1;
logic [RID_WIDTH-1:0] hash_out_2_2;
logic hash_out_valid_filter_2_2;
rule_s_t din_2_2;
rule_s_t din_2_2_r1;
rule_s_t din_2_2_r2;
logic din_valid_2_2;
logic din_valid_2_2_r1;
logic din_valid_2_2_r2;
logic din_almost_full_2_2;
logic [RID_WIDTH-1:0] hash_out_2_3;
logic hash_out_valid_filter_2_3;
rule_s_t din_2_3;
rule_s_t din_2_3_r1;
rule_s_t din_2_3_r2;
logic din_valid_2_3;
logic din_valid_2_3_r1;
logic din_valid_2_3_r2;
logic din_almost_full_2_3;
logic [RID_WIDTH-1:0] hash_out_2_4;
logic hash_out_valid_filter_2_4;
rule_s_t din_2_4;
rule_s_t din_2_4_r1;
rule_s_t din_2_4_r2;
logic din_valid_2_4;
logic din_valid_2_4_r1;
logic din_valid_2_4_r2;
logic din_almost_full_2_4;
logic [RID_WIDTH-1:0] hash_out_2_5;
logic hash_out_valid_filter_2_5;
rule_s_t din_2_5;
rule_s_t din_2_5_r1;
rule_s_t din_2_5_r2;
logic din_valid_2_5;
logic din_valid_2_5_r1;
logic din_valid_2_5_r2;
logic din_almost_full_2_5;
logic [RID_WIDTH-1:0] hash_out_2_6;
logic hash_out_valid_filter_2_6;
rule_s_t din_2_6;
rule_s_t din_2_6_r1;
rule_s_t din_2_6_r2;
logic din_valid_2_6;
logic din_valid_2_6_r1;
logic din_valid_2_6_r2;
logic din_almost_full_2_6;
logic [RID_WIDTH-1:0] hash_out_2_7;
logic hash_out_valid_filter_2_7;
rule_s_t din_2_7;
rule_s_t din_2_7_r1;
rule_s_t din_2_7_r2;
logic din_valid_2_7;
logic din_valid_2_7_r1;
logic din_valid_2_7_r2;
logic din_almost_full_2_7;

rule_s_t din_2_8_r2;
logic din_valid_2_8_r2 = 1'b0;
logic din_almost_full_2_8;
assign din_2_8_r2.data   = 0;
assign din_2_8_r2.last   = 1'b0;
assign din_2_8_r2.bucket = 2;
rule_s_t din_2_9_r2;
logic din_valid_2_9_r2 = 1'b0;
logic din_almost_full_2_9;
assign din_2_9_r2.data   = 0;
assign din_2_9_r2.last   = 1'b0;
assign din_2_9_r2.bucket = 2;
rule_s_t din_2_10_r2;
logic din_valid_2_10_r2 = 1'b0;
logic din_almost_full_2_10;
assign din_2_10_r2.data   = 0;
assign din_2_10_r2.last   = 1'b0;
assign din_2_10_r2.bucket = 2;
rule_s_t din_2_11_r2;
logic din_valid_2_11_r2 = 1'b0;
logic din_almost_full_2_11;
assign din_2_11_r2.data   = 0;
assign din_2_11_r2.last   = 1'b0;
assign din_2_11_r2.bucket = 2;
rule_s_t din_2_12_r2;
logic din_valid_2_12_r2 = 1'b0;
logic din_almost_full_2_12;
assign din_2_12_r2.data   = 0;
assign din_2_12_r2.last   = 1'b0;
assign din_2_12_r2.bucket = 2;
rule_s_t din_2_13_r2;
logic din_valid_2_13_r2 = 1'b0;
logic din_almost_full_2_13;
assign din_2_13_r2.data   = 0;
assign din_2_13_r2.last   = 1'b0;
assign din_2_13_r2.bucket = 2;
rule_s_t din_2_14_r2;
logic din_valid_2_14_r2 = 1'b0;
logic din_almost_full_2_14;
assign din_2_14_r2.data   = 0;
assign din_2_14_r2.last   = 1'b0;
assign din_2_14_r2.bucket = 2;
rule_s_t din_2_15_r2;
logic din_valid_2_15_r2 = 1'b0;
logic din_almost_full_2_15;
assign din_2_15_r2.data   = 0;
assign din_2_15_r2.last   = 1'b0;
assign din_2_15_r2.bucket = 2;
rule_s_t din_2_16_r2;
logic din_valid_2_16_r2 = 1'b0;
logic din_almost_full_2_16;
assign din_2_16_r2.data   = 0;
assign din_2_16_r2.last   = 1'b0;
assign din_2_16_r2.bucket = 2;
rule_s_t din_2_17_r2;
logic din_valid_2_17_r2 = 1'b0;
logic din_almost_full_2_17;
assign din_2_17_r2.data   = 0;
assign din_2_17_r2.last   = 1'b0;
assign din_2_17_r2.bucket = 2;
rule_s_t din_2_18_r2;
logic din_valid_2_18_r2 = 1'b0;
logic din_almost_full_2_18;
assign din_2_18_r2.data   = 0;
assign din_2_18_r2.last   = 1'b0;
assign din_2_18_r2.bucket = 2;
rule_s_t din_2_19_r2;
logic din_valid_2_19_r2 = 1'b0;
logic din_almost_full_2_19;
assign din_2_19_r2.data   = 0;
assign din_2_19_r2.last   = 1'b0;
assign din_2_19_r2.bucket = 2;
rule_s_t din_2_20_r2;
logic din_valid_2_20_r2 = 1'b0;
logic din_almost_full_2_20;
assign din_2_20_r2.data   = 0;
assign din_2_20_r2.last   = 1'b0;
assign din_2_20_r2.bucket = 2;
rule_s_t din_2_21_r2;
logic din_valid_2_21_r2 = 1'b0;
logic din_almost_full_2_21;
assign din_2_21_r2.data   = 0;
assign din_2_21_r2.last   = 1'b0;
assign din_2_21_r2.bucket = 2;
rule_s_t din_2_22_r2;
logic din_valid_2_22_r2 = 1'b0;
logic din_almost_full_2_22;
assign din_2_22_r2.data   = 0;
assign din_2_22_r2.last   = 1'b0;
assign din_2_22_r2.bucket = 2;
rule_s_t din_2_23_r2;
logic din_valid_2_23_r2 = 1'b0;
logic din_almost_full_2_23;
assign din_2_23_r2.data   = 0;
assign din_2_23_r2.last   = 1'b0;
assign din_2_23_r2.bucket = 2;
rule_s_t din_2_24_r2;
logic din_valid_2_24_r2 = 1'b0;
logic din_almost_full_2_24;
assign din_2_24_r2.data   = 0;
assign din_2_24_r2.last   = 1'b0;
assign din_2_24_r2.bucket = 2;
rule_s_t din_2_25_r2;
logic din_valid_2_25_r2 = 1'b0;
logic din_almost_full_2_25;
assign din_2_25_r2.data   = 0;
assign din_2_25_r2.last   = 1'b0;
assign din_2_25_r2.bucket = 2;
rule_s_t din_2_26_r2;
logic din_valid_2_26_r2 = 1'b0;
logic din_almost_full_2_26;
assign din_2_26_r2.data   = 0;
assign din_2_26_r2.last   = 1'b0;
assign din_2_26_r2.bucket = 2;
rule_s_t din_2_27_r2;
logic din_valid_2_27_r2 = 1'b0;
logic din_almost_full_2_27;
assign din_2_27_r2.data   = 0;
assign din_2_27_r2.last   = 1'b0;
assign din_2_27_r2.bucket = 2;
rule_s_t din_2_28_r2;
logic din_valid_2_28_r2 = 1'b0;
logic din_almost_full_2_28;
assign din_2_28_r2.data   = 0;
assign din_2_28_r2.last   = 1'b0;
assign din_2_28_r2.bucket = 2;
rule_s_t din_2_29_r2;
logic din_valid_2_29_r2 = 1'b0;
logic din_almost_full_2_29;
assign din_2_29_r2.data   = 0;
assign din_2_29_r2.last   = 1'b0;
assign din_2_29_r2.bucket = 2;
rule_s_t din_2_30_r2;
logic din_valid_2_30_r2 = 1'b0;
logic din_almost_full_2_30;
assign din_2_30_r2.data   = 0;
assign din_2_30_r2.last   = 1'b0;
assign din_2_30_r2.bucket = 2;
rule_s_t din_2_31_r2;
logic din_valid_2_31_r2 = 1'b0;
logic din_almost_full_2_31;
assign din_2_31_r2.data   = 0;
assign din_2_31_r2.last   = 1'b0;
assign din_2_31_r2.bucket = 2;

logic [RID_WIDTH-1:0] hash_out_3_0;
logic hash_out_valid_filter_3_0;
rule_s_t din_3_0;
rule_s_t din_3_0_r1;
rule_s_t din_3_0_r2;
logic din_valid_3_0;
logic din_valid_3_0_r1;
logic din_valid_3_0_r2;
logic din_almost_full_3_0;
logic [RID_WIDTH-1:0] hash_out_3_1;
logic hash_out_valid_filter_3_1;
rule_s_t din_3_1;
rule_s_t din_3_1_r1;
rule_s_t din_3_1_r2;
logic din_valid_3_1;
logic din_valid_3_1_r1;
logic din_valid_3_1_r2;
logic din_almost_full_3_1;
logic [RID_WIDTH-1:0] hash_out_3_2;
logic hash_out_valid_filter_3_2;
rule_s_t din_3_2;
rule_s_t din_3_2_r1;
rule_s_t din_3_2_r2;
logic din_valid_3_2;
logic din_valid_3_2_r1;
logic din_valid_3_2_r2;
logic din_almost_full_3_2;
logic [RID_WIDTH-1:0] hash_out_3_3;
logic hash_out_valid_filter_3_3;
rule_s_t din_3_3;
rule_s_t din_3_3_r1;
rule_s_t din_3_3_r2;
logic din_valid_3_3;
logic din_valid_3_3_r1;
logic din_valid_3_3_r2;
logic din_almost_full_3_3;
logic [RID_WIDTH-1:0] hash_out_3_4;
logic hash_out_valid_filter_3_4;
rule_s_t din_3_4;
rule_s_t din_3_4_r1;
rule_s_t din_3_4_r2;
logic din_valid_3_4;
logic din_valid_3_4_r1;
logic din_valid_3_4_r2;
logic din_almost_full_3_4;
logic [RID_WIDTH-1:0] hash_out_3_5;
logic hash_out_valid_filter_3_5;
rule_s_t din_3_5;
rule_s_t din_3_5_r1;
rule_s_t din_3_5_r2;
logic din_valid_3_5;
logic din_valid_3_5_r1;
logic din_valid_3_5_r2;
logic din_almost_full_3_5;
logic [RID_WIDTH-1:0] hash_out_3_6;
logic hash_out_valid_filter_3_6;
rule_s_t din_3_6;
rule_s_t din_3_6_r1;
rule_s_t din_3_6_r2;
logic din_valid_3_6;
logic din_valid_3_6_r1;
logic din_valid_3_6_r2;
logic din_almost_full_3_6;
logic [RID_WIDTH-1:0] hash_out_3_7;
logic hash_out_valid_filter_3_7;
rule_s_t din_3_7;
rule_s_t din_3_7_r1;
rule_s_t din_3_7_r2;
logic din_valid_3_7;
logic din_valid_3_7_r1;
logic din_valid_3_7_r2;
logic din_almost_full_3_7;

rule_s_t din_3_8_r2;
logic din_valid_3_8_r2 = 1'b0;
logic din_almost_full_3_8;
assign din_3_8_r2.data   = 0;
assign din_3_8_r2.last   = 1'b0;
assign din_3_8_r2.bucket = 3;
rule_s_t din_3_9_r2;
logic din_valid_3_9_r2 = 1'b0;
logic din_almost_full_3_9;
assign din_3_9_r2.data   = 0;
assign din_3_9_r2.last   = 1'b0;
assign din_3_9_r2.bucket = 3;
rule_s_t din_3_10_r2;
logic din_valid_3_10_r2 = 1'b0;
logic din_almost_full_3_10;
assign din_3_10_r2.data   = 0;
assign din_3_10_r2.last   = 1'b0;
assign din_3_10_r2.bucket = 3;
rule_s_t din_3_11_r2;
logic din_valid_3_11_r2 = 1'b0;
logic din_almost_full_3_11;
assign din_3_11_r2.data   = 0;
assign din_3_11_r2.last   = 1'b0;
assign din_3_11_r2.bucket = 3;
rule_s_t din_3_12_r2;
logic din_valid_3_12_r2 = 1'b0;
logic din_almost_full_3_12;
assign din_3_12_r2.data   = 0;
assign din_3_12_r2.last   = 1'b0;
assign din_3_12_r2.bucket = 3;
rule_s_t din_3_13_r2;
logic din_valid_3_13_r2 = 1'b0;
logic din_almost_full_3_13;
assign din_3_13_r2.data   = 0;
assign din_3_13_r2.last   = 1'b0;
assign din_3_13_r2.bucket = 3;
rule_s_t din_3_14_r2;
logic din_valid_3_14_r2 = 1'b0;
logic din_almost_full_3_14;
assign din_3_14_r2.data   = 0;
assign din_3_14_r2.last   = 1'b0;
assign din_3_14_r2.bucket = 3;
rule_s_t din_3_15_r2;
logic din_valid_3_15_r2 = 1'b0;
logic din_almost_full_3_15;
assign din_3_15_r2.data   = 0;
assign din_3_15_r2.last   = 1'b0;
assign din_3_15_r2.bucket = 3;
rule_s_t din_3_16_r2;
logic din_valid_3_16_r2 = 1'b0;
logic din_almost_full_3_16;
assign din_3_16_r2.data   = 0;
assign din_3_16_r2.last   = 1'b0;
assign din_3_16_r2.bucket = 3;
rule_s_t din_3_17_r2;
logic din_valid_3_17_r2 = 1'b0;
logic din_almost_full_3_17;
assign din_3_17_r2.data   = 0;
assign din_3_17_r2.last   = 1'b0;
assign din_3_17_r2.bucket = 3;
rule_s_t din_3_18_r2;
logic din_valid_3_18_r2 = 1'b0;
logic din_almost_full_3_18;
assign din_3_18_r2.data   = 0;
assign din_3_18_r2.last   = 1'b0;
assign din_3_18_r2.bucket = 3;
rule_s_t din_3_19_r2;
logic din_valid_3_19_r2 = 1'b0;
logic din_almost_full_3_19;
assign din_3_19_r2.data   = 0;
assign din_3_19_r2.last   = 1'b0;
assign din_3_19_r2.bucket = 3;
rule_s_t din_3_20_r2;
logic din_valid_3_20_r2 = 1'b0;
logic din_almost_full_3_20;
assign din_3_20_r2.data   = 0;
assign din_3_20_r2.last   = 1'b0;
assign din_3_20_r2.bucket = 3;
rule_s_t din_3_21_r2;
logic din_valid_3_21_r2 = 1'b0;
logic din_almost_full_3_21;
assign din_3_21_r2.data   = 0;
assign din_3_21_r2.last   = 1'b0;
assign din_3_21_r2.bucket = 3;
rule_s_t din_3_22_r2;
logic din_valid_3_22_r2 = 1'b0;
logic din_almost_full_3_22;
assign din_3_22_r2.data   = 0;
assign din_3_22_r2.last   = 1'b0;
assign din_3_22_r2.bucket = 3;
rule_s_t din_3_23_r2;
logic din_valid_3_23_r2 = 1'b0;
logic din_almost_full_3_23;
assign din_3_23_r2.data   = 0;
assign din_3_23_r2.last   = 1'b0;
assign din_3_23_r2.bucket = 3;
rule_s_t din_3_24_r2;
logic din_valid_3_24_r2 = 1'b0;
logic din_almost_full_3_24;
assign din_3_24_r2.data   = 0;
assign din_3_24_r2.last   = 1'b0;
assign din_3_24_r2.bucket = 3;
rule_s_t din_3_25_r2;
logic din_valid_3_25_r2 = 1'b0;
logic din_almost_full_3_25;
assign din_3_25_r2.data   = 0;
assign din_3_25_r2.last   = 1'b0;
assign din_3_25_r2.bucket = 3;
rule_s_t din_3_26_r2;
logic din_valid_3_26_r2 = 1'b0;
logic din_almost_full_3_26;
assign din_3_26_r2.data   = 0;
assign din_3_26_r2.last   = 1'b0;
assign din_3_26_r2.bucket = 3;
rule_s_t din_3_27_r2;
logic din_valid_3_27_r2 = 1'b0;
logic din_almost_full_3_27;
assign din_3_27_r2.data   = 0;
assign din_3_27_r2.last   = 1'b0;
assign din_3_27_r2.bucket = 3;
rule_s_t din_3_28_r2;
logic din_valid_3_28_r2 = 1'b0;
logic din_almost_full_3_28;
assign din_3_28_r2.data   = 0;
assign din_3_28_r2.last   = 1'b0;
assign din_3_28_r2.bucket = 3;
rule_s_t din_3_29_r2;
logic din_valid_3_29_r2 = 1'b0;
logic din_almost_full_3_29;
assign din_3_29_r2.data   = 0;
assign din_3_29_r2.last   = 1'b0;
assign din_3_29_r2.bucket = 3;
rule_s_t din_3_30_r2;
logic din_valid_3_30_r2 = 1'b0;
logic din_almost_full_3_30;
assign din_3_30_r2.data   = 0;
assign din_3_30_r2.last   = 1'b0;
assign din_3_30_r2.bucket = 3;
rule_s_t din_3_31_r2;
logic din_valid_3_31_r2 = 1'b0;
logic din_almost_full_3_31;
assign din_3_31_r2.data   = 0;
assign din_3_31_r2.last   = 1'b0;
assign din_3_31_r2.bucket = 3;

logic [RID_WIDTH-1:0] hash_out_4_0;
logic hash_out_valid_filter_4_0;
rule_s_t din_4_0;
rule_s_t din_4_0_r1;
rule_s_t din_4_0_r2;
logic din_valid_4_0;
logic din_valid_4_0_r1;
logic din_valid_4_0_r2;
logic din_almost_full_4_0;
logic [RID_WIDTH-1:0] hash_out_4_1;
logic hash_out_valid_filter_4_1;
rule_s_t din_4_1;
rule_s_t din_4_1_r1;
rule_s_t din_4_1_r2;
logic din_valid_4_1;
logic din_valid_4_1_r1;
logic din_valid_4_1_r2;
logic din_almost_full_4_1;
logic [RID_WIDTH-1:0] hash_out_4_2;
logic hash_out_valid_filter_4_2;
rule_s_t din_4_2;
rule_s_t din_4_2_r1;
rule_s_t din_4_2_r2;
logic din_valid_4_2;
logic din_valid_4_2_r1;
logic din_valid_4_2_r2;
logic din_almost_full_4_2;
logic [RID_WIDTH-1:0] hash_out_4_3;
logic hash_out_valid_filter_4_3;
rule_s_t din_4_3;
rule_s_t din_4_3_r1;
rule_s_t din_4_3_r2;
logic din_valid_4_3;
logic din_valid_4_3_r1;
logic din_valid_4_3_r2;
logic din_almost_full_4_3;
logic [RID_WIDTH-1:0] hash_out_4_4;
logic hash_out_valid_filter_4_4;
rule_s_t din_4_4;
rule_s_t din_4_4_r1;
rule_s_t din_4_4_r2;
logic din_valid_4_4;
logic din_valid_4_4_r1;
logic din_valid_4_4_r2;
logic din_almost_full_4_4;
logic [RID_WIDTH-1:0] hash_out_4_5;
logic hash_out_valid_filter_4_5;
rule_s_t din_4_5;
rule_s_t din_4_5_r1;
rule_s_t din_4_5_r2;
logic din_valid_4_5;
logic din_valid_4_5_r1;
logic din_valid_4_5_r2;
logic din_almost_full_4_5;
logic [RID_WIDTH-1:0] hash_out_4_6;
logic hash_out_valid_filter_4_6;
rule_s_t din_4_6;
rule_s_t din_4_6_r1;
rule_s_t din_4_6_r2;
logic din_valid_4_6;
logic din_valid_4_6_r1;
logic din_valid_4_6_r2;
logic din_almost_full_4_6;
logic [RID_WIDTH-1:0] hash_out_4_7;
logic hash_out_valid_filter_4_7;
rule_s_t din_4_7;
rule_s_t din_4_7_r1;
rule_s_t din_4_7_r2;
logic din_valid_4_7;
logic din_valid_4_7_r1;
logic din_valid_4_7_r2;
logic din_almost_full_4_7;

rule_s_t din_4_8_r2;
logic din_valid_4_8_r2 = 1'b0;
logic din_almost_full_4_8;
assign din_4_8_r2.data   = 0;
assign din_4_8_r2.last   = 1'b0;
assign din_4_8_r2.bucket = 4;
rule_s_t din_4_9_r2;
logic din_valid_4_9_r2 = 1'b0;
logic din_almost_full_4_9;
assign din_4_9_r2.data   = 0;
assign din_4_9_r2.last   = 1'b0;
assign din_4_9_r2.bucket = 4;
rule_s_t din_4_10_r2;
logic din_valid_4_10_r2 = 1'b0;
logic din_almost_full_4_10;
assign din_4_10_r2.data   = 0;
assign din_4_10_r2.last   = 1'b0;
assign din_4_10_r2.bucket = 4;
rule_s_t din_4_11_r2;
logic din_valid_4_11_r2 = 1'b0;
logic din_almost_full_4_11;
assign din_4_11_r2.data   = 0;
assign din_4_11_r2.last   = 1'b0;
assign din_4_11_r2.bucket = 4;
rule_s_t din_4_12_r2;
logic din_valid_4_12_r2 = 1'b0;
logic din_almost_full_4_12;
assign din_4_12_r2.data   = 0;
assign din_4_12_r2.last   = 1'b0;
assign din_4_12_r2.bucket = 4;
rule_s_t din_4_13_r2;
logic din_valid_4_13_r2 = 1'b0;
logic din_almost_full_4_13;
assign din_4_13_r2.data   = 0;
assign din_4_13_r2.last   = 1'b0;
assign din_4_13_r2.bucket = 4;
rule_s_t din_4_14_r2;
logic din_valid_4_14_r2 = 1'b0;
logic din_almost_full_4_14;
assign din_4_14_r2.data   = 0;
assign din_4_14_r2.last   = 1'b0;
assign din_4_14_r2.bucket = 4;
rule_s_t din_4_15_r2;
logic din_valid_4_15_r2 = 1'b0;
logic din_almost_full_4_15;
assign din_4_15_r2.data   = 0;
assign din_4_15_r2.last   = 1'b0;
assign din_4_15_r2.bucket = 4;
rule_s_t din_4_16_r2;
logic din_valid_4_16_r2 = 1'b0;
logic din_almost_full_4_16;
assign din_4_16_r2.data   = 0;
assign din_4_16_r2.last   = 1'b0;
assign din_4_16_r2.bucket = 4;
rule_s_t din_4_17_r2;
logic din_valid_4_17_r2 = 1'b0;
logic din_almost_full_4_17;
assign din_4_17_r2.data   = 0;
assign din_4_17_r2.last   = 1'b0;
assign din_4_17_r2.bucket = 4;
rule_s_t din_4_18_r2;
logic din_valid_4_18_r2 = 1'b0;
logic din_almost_full_4_18;
assign din_4_18_r2.data   = 0;
assign din_4_18_r2.last   = 1'b0;
assign din_4_18_r2.bucket = 4;
rule_s_t din_4_19_r2;
logic din_valid_4_19_r2 = 1'b0;
logic din_almost_full_4_19;
assign din_4_19_r2.data   = 0;
assign din_4_19_r2.last   = 1'b0;
assign din_4_19_r2.bucket = 4;
rule_s_t din_4_20_r2;
logic din_valid_4_20_r2 = 1'b0;
logic din_almost_full_4_20;
assign din_4_20_r2.data   = 0;
assign din_4_20_r2.last   = 1'b0;
assign din_4_20_r2.bucket = 4;
rule_s_t din_4_21_r2;
logic din_valid_4_21_r2 = 1'b0;
logic din_almost_full_4_21;
assign din_4_21_r2.data   = 0;
assign din_4_21_r2.last   = 1'b0;
assign din_4_21_r2.bucket = 4;
rule_s_t din_4_22_r2;
logic din_valid_4_22_r2 = 1'b0;
logic din_almost_full_4_22;
assign din_4_22_r2.data   = 0;
assign din_4_22_r2.last   = 1'b0;
assign din_4_22_r2.bucket = 4;
rule_s_t din_4_23_r2;
logic din_valid_4_23_r2 = 1'b0;
logic din_almost_full_4_23;
assign din_4_23_r2.data   = 0;
assign din_4_23_r2.last   = 1'b0;
assign din_4_23_r2.bucket = 4;
rule_s_t din_4_24_r2;
logic din_valid_4_24_r2 = 1'b0;
logic din_almost_full_4_24;
assign din_4_24_r2.data   = 0;
assign din_4_24_r2.last   = 1'b0;
assign din_4_24_r2.bucket = 4;
rule_s_t din_4_25_r2;
logic din_valid_4_25_r2 = 1'b0;
logic din_almost_full_4_25;
assign din_4_25_r2.data   = 0;
assign din_4_25_r2.last   = 1'b0;
assign din_4_25_r2.bucket = 4;
rule_s_t din_4_26_r2;
logic din_valid_4_26_r2 = 1'b0;
logic din_almost_full_4_26;
assign din_4_26_r2.data   = 0;
assign din_4_26_r2.last   = 1'b0;
assign din_4_26_r2.bucket = 4;
rule_s_t din_4_27_r2;
logic din_valid_4_27_r2 = 1'b0;
logic din_almost_full_4_27;
assign din_4_27_r2.data   = 0;
assign din_4_27_r2.last   = 1'b0;
assign din_4_27_r2.bucket = 4;
rule_s_t din_4_28_r2;
logic din_valid_4_28_r2 = 1'b0;
logic din_almost_full_4_28;
assign din_4_28_r2.data   = 0;
assign din_4_28_r2.last   = 1'b0;
assign din_4_28_r2.bucket = 4;
rule_s_t din_4_29_r2;
logic din_valid_4_29_r2 = 1'b0;
logic din_almost_full_4_29;
assign din_4_29_r2.data   = 0;
assign din_4_29_r2.last   = 1'b0;
assign din_4_29_r2.bucket = 4;
rule_s_t din_4_30_r2;
logic din_valid_4_30_r2 = 1'b0;
logic din_almost_full_4_30;
assign din_4_30_r2.data   = 0;
assign din_4_30_r2.last   = 1'b0;
assign din_4_30_r2.bucket = 4;
rule_s_t din_4_31_r2;
logic din_valid_4_31_r2 = 1'b0;
logic din_almost_full_4_31;
assign din_4_31_r2.data   = 0;
assign din_4_31_r2.last   = 1'b0;
assign din_4_31_r2.bucket = 4;

logic [RID_WIDTH-1:0] hash_out_5_0;
logic hash_out_valid_filter_5_0;
rule_s_t din_5_0;
rule_s_t din_5_0_r1;
rule_s_t din_5_0_r2;
logic din_valid_5_0;
logic din_valid_5_0_r1;
logic din_valid_5_0_r2;
logic din_almost_full_5_0;
logic [RID_WIDTH-1:0] hash_out_5_1;
logic hash_out_valid_filter_5_1;
rule_s_t din_5_1;
rule_s_t din_5_1_r1;
rule_s_t din_5_1_r2;
logic din_valid_5_1;
logic din_valid_5_1_r1;
logic din_valid_5_1_r2;
logic din_almost_full_5_1;
logic [RID_WIDTH-1:0] hash_out_5_2;
logic hash_out_valid_filter_5_2;
rule_s_t din_5_2;
rule_s_t din_5_2_r1;
rule_s_t din_5_2_r2;
logic din_valid_5_2;
logic din_valid_5_2_r1;
logic din_valid_5_2_r2;
logic din_almost_full_5_2;
logic [RID_WIDTH-1:0] hash_out_5_3;
logic hash_out_valid_filter_5_3;
rule_s_t din_5_3;
rule_s_t din_5_3_r1;
rule_s_t din_5_3_r2;
logic din_valid_5_3;
logic din_valid_5_3_r1;
logic din_valid_5_3_r2;
logic din_almost_full_5_3;
logic [RID_WIDTH-1:0] hash_out_5_4;
logic hash_out_valid_filter_5_4;
rule_s_t din_5_4;
rule_s_t din_5_4_r1;
rule_s_t din_5_4_r2;
logic din_valid_5_4;
logic din_valid_5_4_r1;
logic din_valid_5_4_r2;
logic din_almost_full_5_4;
logic [RID_WIDTH-1:0] hash_out_5_5;
logic hash_out_valid_filter_5_5;
rule_s_t din_5_5;
rule_s_t din_5_5_r1;
rule_s_t din_5_5_r2;
logic din_valid_5_5;
logic din_valid_5_5_r1;
logic din_valid_5_5_r2;
logic din_almost_full_5_5;
logic [RID_WIDTH-1:0] hash_out_5_6;
logic hash_out_valid_filter_5_6;
rule_s_t din_5_6;
rule_s_t din_5_6_r1;
rule_s_t din_5_6_r2;
logic din_valid_5_6;
logic din_valid_5_6_r1;
logic din_valid_5_6_r2;
logic din_almost_full_5_6;
logic [RID_WIDTH-1:0] hash_out_5_7;
logic hash_out_valid_filter_5_7;
rule_s_t din_5_7;
rule_s_t din_5_7_r1;
rule_s_t din_5_7_r2;
logic din_valid_5_7;
logic din_valid_5_7_r1;
logic din_valid_5_7_r2;
logic din_almost_full_5_7;

rule_s_t din_5_8_r2;
logic din_valid_5_8_r2 = 1'b0;
logic din_almost_full_5_8;
assign din_5_8_r2.data   = 0;
assign din_5_8_r2.last   = 1'b0;
assign din_5_8_r2.bucket = 5;
rule_s_t din_5_9_r2;
logic din_valid_5_9_r2 = 1'b0;
logic din_almost_full_5_9;
assign din_5_9_r2.data   = 0;
assign din_5_9_r2.last   = 1'b0;
assign din_5_9_r2.bucket = 5;
rule_s_t din_5_10_r2;
logic din_valid_5_10_r2 = 1'b0;
logic din_almost_full_5_10;
assign din_5_10_r2.data   = 0;
assign din_5_10_r2.last   = 1'b0;
assign din_5_10_r2.bucket = 5;
rule_s_t din_5_11_r2;
logic din_valid_5_11_r2 = 1'b0;
logic din_almost_full_5_11;
assign din_5_11_r2.data   = 0;
assign din_5_11_r2.last   = 1'b0;
assign din_5_11_r2.bucket = 5;
rule_s_t din_5_12_r2;
logic din_valid_5_12_r2 = 1'b0;
logic din_almost_full_5_12;
assign din_5_12_r2.data   = 0;
assign din_5_12_r2.last   = 1'b0;
assign din_5_12_r2.bucket = 5;
rule_s_t din_5_13_r2;
logic din_valid_5_13_r2 = 1'b0;
logic din_almost_full_5_13;
assign din_5_13_r2.data   = 0;
assign din_5_13_r2.last   = 1'b0;
assign din_5_13_r2.bucket = 5;
rule_s_t din_5_14_r2;
logic din_valid_5_14_r2 = 1'b0;
logic din_almost_full_5_14;
assign din_5_14_r2.data   = 0;
assign din_5_14_r2.last   = 1'b0;
assign din_5_14_r2.bucket = 5;
rule_s_t din_5_15_r2;
logic din_valid_5_15_r2 = 1'b0;
logic din_almost_full_5_15;
assign din_5_15_r2.data   = 0;
assign din_5_15_r2.last   = 1'b0;
assign din_5_15_r2.bucket = 5;
rule_s_t din_5_16_r2;
logic din_valid_5_16_r2 = 1'b0;
logic din_almost_full_5_16;
assign din_5_16_r2.data   = 0;
assign din_5_16_r2.last   = 1'b0;
assign din_5_16_r2.bucket = 5;
rule_s_t din_5_17_r2;
logic din_valid_5_17_r2 = 1'b0;
logic din_almost_full_5_17;
assign din_5_17_r2.data   = 0;
assign din_5_17_r2.last   = 1'b0;
assign din_5_17_r2.bucket = 5;
rule_s_t din_5_18_r2;
logic din_valid_5_18_r2 = 1'b0;
logic din_almost_full_5_18;
assign din_5_18_r2.data   = 0;
assign din_5_18_r2.last   = 1'b0;
assign din_5_18_r2.bucket = 5;
rule_s_t din_5_19_r2;
logic din_valid_5_19_r2 = 1'b0;
logic din_almost_full_5_19;
assign din_5_19_r2.data   = 0;
assign din_5_19_r2.last   = 1'b0;
assign din_5_19_r2.bucket = 5;
rule_s_t din_5_20_r2;
logic din_valid_5_20_r2 = 1'b0;
logic din_almost_full_5_20;
assign din_5_20_r2.data   = 0;
assign din_5_20_r2.last   = 1'b0;
assign din_5_20_r2.bucket = 5;
rule_s_t din_5_21_r2;
logic din_valid_5_21_r2 = 1'b0;
logic din_almost_full_5_21;
assign din_5_21_r2.data   = 0;
assign din_5_21_r2.last   = 1'b0;
assign din_5_21_r2.bucket = 5;
rule_s_t din_5_22_r2;
logic din_valid_5_22_r2 = 1'b0;
logic din_almost_full_5_22;
assign din_5_22_r2.data   = 0;
assign din_5_22_r2.last   = 1'b0;
assign din_5_22_r2.bucket = 5;
rule_s_t din_5_23_r2;
logic din_valid_5_23_r2 = 1'b0;
logic din_almost_full_5_23;
assign din_5_23_r2.data   = 0;
assign din_5_23_r2.last   = 1'b0;
assign din_5_23_r2.bucket = 5;
rule_s_t din_5_24_r2;
logic din_valid_5_24_r2 = 1'b0;
logic din_almost_full_5_24;
assign din_5_24_r2.data   = 0;
assign din_5_24_r2.last   = 1'b0;
assign din_5_24_r2.bucket = 5;
rule_s_t din_5_25_r2;
logic din_valid_5_25_r2 = 1'b0;
logic din_almost_full_5_25;
assign din_5_25_r2.data   = 0;
assign din_5_25_r2.last   = 1'b0;
assign din_5_25_r2.bucket = 5;
rule_s_t din_5_26_r2;
logic din_valid_5_26_r2 = 1'b0;
logic din_almost_full_5_26;
assign din_5_26_r2.data   = 0;
assign din_5_26_r2.last   = 1'b0;
assign din_5_26_r2.bucket = 5;
rule_s_t din_5_27_r2;
logic din_valid_5_27_r2 = 1'b0;
logic din_almost_full_5_27;
assign din_5_27_r2.data   = 0;
assign din_5_27_r2.last   = 1'b0;
assign din_5_27_r2.bucket = 5;
rule_s_t din_5_28_r2;
logic din_valid_5_28_r2 = 1'b0;
logic din_almost_full_5_28;
assign din_5_28_r2.data   = 0;
assign din_5_28_r2.last   = 1'b0;
assign din_5_28_r2.bucket = 5;
rule_s_t din_5_29_r2;
logic din_valid_5_29_r2 = 1'b0;
logic din_almost_full_5_29;
assign din_5_29_r2.data   = 0;
assign din_5_29_r2.last   = 1'b0;
assign din_5_29_r2.bucket = 5;
rule_s_t din_5_30_r2;
logic din_valid_5_30_r2 = 1'b0;
logic din_almost_full_5_30;
assign din_5_30_r2.data   = 0;
assign din_5_30_r2.last   = 1'b0;
assign din_5_30_r2.bucket = 5;
rule_s_t din_5_31_r2;
logic din_valid_5_31_r2 = 1'b0;
logic din_almost_full_5_31;
assign din_5_31_r2.data   = 0;
assign din_5_31_r2.last   = 1'b0;
assign din_5_31_r2.bucket = 5;

logic [RID_WIDTH-1:0] hash_out_6_0;
logic hash_out_valid_filter_6_0;
rule_s_t din_6_0;
rule_s_t din_6_0_r1;
rule_s_t din_6_0_r2;
logic din_valid_6_0;
logic din_valid_6_0_r1;
logic din_valid_6_0_r2;
logic din_almost_full_6_0;
logic [RID_WIDTH-1:0] hash_out_6_1;
logic hash_out_valid_filter_6_1;
rule_s_t din_6_1;
rule_s_t din_6_1_r1;
rule_s_t din_6_1_r2;
logic din_valid_6_1;
logic din_valid_6_1_r1;
logic din_valid_6_1_r2;
logic din_almost_full_6_1;
logic [RID_WIDTH-1:0] hash_out_6_2;
logic hash_out_valid_filter_6_2;
rule_s_t din_6_2;
rule_s_t din_6_2_r1;
rule_s_t din_6_2_r2;
logic din_valid_6_2;
logic din_valid_6_2_r1;
logic din_valid_6_2_r2;
logic din_almost_full_6_2;
logic [RID_WIDTH-1:0] hash_out_6_3;
logic hash_out_valid_filter_6_3;
rule_s_t din_6_3;
rule_s_t din_6_3_r1;
rule_s_t din_6_3_r2;
logic din_valid_6_3;
logic din_valid_6_3_r1;
logic din_valid_6_3_r2;
logic din_almost_full_6_3;
logic [RID_WIDTH-1:0] hash_out_6_4;
logic hash_out_valid_filter_6_4;
rule_s_t din_6_4;
rule_s_t din_6_4_r1;
rule_s_t din_6_4_r2;
logic din_valid_6_4;
logic din_valid_6_4_r1;
logic din_valid_6_4_r2;
logic din_almost_full_6_4;
logic [RID_WIDTH-1:0] hash_out_6_5;
logic hash_out_valid_filter_6_5;
rule_s_t din_6_5;
rule_s_t din_6_5_r1;
rule_s_t din_6_5_r2;
logic din_valid_6_5;
logic din_valid_6_5_r1;
logic din_valid_6_5_r2;
logic din_almost_full_6_5;
logic [RID_WIDTH-1:0] hash_out_6_6;
logic hash_out_valid_filter_6_6;
rule_s_t din_6_6;
rule_s_t din_6_6_r1;
rule_s_t din_6_6_r2;
logic din_valid_6_6;
logic din_valid_6_6_r1;
logic din_valid_6_6_r2;
logic din_almost_full_6_6;
logic [RID_WIDTH-1:0] hash_out_6_7;
logic hash_out_valid_filter_6_7;
rule_s_t din_6_7;
rule_s_t din_6_7_r1;
rule_s_t din_6_7_r2;
logic din_valid_6_7;
logic din_valid_6_7_r1;
logic din_valid_6_7_r2;
logic din_almost_full_6_7;

rule_s_t din_6_8_r2;
logic din_valid_6_8_r2 = 1'b0;
logic din_almost_full_6_8;
assign din_6_8_r2.data   = 0;
assign din_6_8_r2.last   = 1'b0;
assign din_6_8_r2.bucket = 6;
rule_s_t din_6_9_r2;
logic din_valid_6_9_r2 = 1'b0;
logic din_almost_full_6_9;
assign din_6_9_r2.data   = 0;
assign din_6_9_r2.last   = 1'b0;
assign din_6_9_r2.bucket = 6;
rule_s_t din_6_10_r2;
logic din_valid_6_10_r2 = 1'b0;
logic din_almost_full_6_10;
assign din_6_10_r2.data   = 0;
assign din_6_10_r2.last   = 1'b0;
assign din_6_10_r2.bucket = 6;
rule_s_t din_6_11_r2;
logic din_valid_6_11_r2 = 1'b0;
logic din_almost_full_6_11;
assign din_6_11_r2.data   = 0;
assign din_6_11_r2.last   = 1'b0;
assign din_6_11_r2.bucket = 6;
rule_s_t din_6_12_r2;
logic din_valid_6_12_r2 = 1'b0;
logic din_almost_full_6_12;
assign din_6_12_r2.data   = 0;
assign din_6_12_r2.last   = 1'b0;
assign din_6_12_r2.bucket = 6;
rule_s_t din_6_13_r2;
logic din_valid_6_13_r2 = 1'b0;
logic din_almost_full_6_13;
assign din_6_13_r2.data   = 0;
assign din_6_13_r2.last   = 1'b0;
assign din_6_13_r2.bucket = 6;
rule_s_t din_6_14_r2;
logic din_valid_6_14_r2 = 1'b0;
logic din_almost_full_6_14;
assign din_6_14_r2.data   = 0;
assign din_6_14_r2.last   = 1'b0;
assign din_6_14_r2.bucket = 6;
rule_s_t din_6_15_r2;
logic din_valid_6_15_r2 = 1'b0;
logic din_almost_full_6_15;
assign din_6_15_r2.data   = 0;
assign din_6_15_r2.last   = 1'b0;
assign din_6_15_r2.bucket = 6;
rule_s_t din_6_16_r2;
logic din_valid_6_16_r2 = 1'b0;
logic din_almost_full_6_16;
assign din_6_16_r2.data   = 0;
assign din_6_16_r2.last   = 1'b0;
assign din_6_16_r2.bucket = 6;
rule_s_t din_6_17_r2;
logic din_valid_6_17_r2 = 1'b0;
logic din_almost_full_6_17;
assign din_6_17_r2.data   = 0;
assign din_6_17_r2.last   = 1'b0;
assign din_6_17_r2.bucket = 6;
rule_s_t din_6_18_r2;
logic din_valid_6_18_r2 = 1'b0;
logic din_almost_full_6_18;
assign din_6_18_r2.data   = 0;
assign din_6_18_r2.last   = 1'b0;
assign din_6_18_r2.bucket = 6;
rule_s_t din_6_19_r2;
logic din_valid_6_19_r2 = 1'b0;
logic din_almost_full_6_19;
assign din_6_19_r2.data   = 0;
assign din_6_19_r2.last   = 1'b0;
assign din_6_19_r2.bucket = 6;
rule_s_t din_6_20_r2;
logic din_valid_6_20_r2 = 1'b0;
logic din_almost_full_6_20;
assign din_6_20_r2.data   = 0;
assign din_6_20_r2.last   = 1'b0;
assign din_6_20_r2.bucket = 6;
rule_s_t din_6_21_r2;
logic din_valid_6_21_r2 = 1'b0;
logic din_almost_full_6_21;
assign din_6_21_r2.data   = 0;
assign din_6_21_r2.last   = 1'b0;
assign din_6_21_r2.bucket = 6;
rule_s_t din_6_22_r2;
logic din_valid_6_22_r2 = 1'b0;
logic din_almost_full_6_22;
assign din_6_22_r2.data   = 0;
assign din_6_22_r2.last   = 1'b0;
assign din_6_22_r2.bucket = 6;
rule_s_t din_6_23_r2;
logic din_valid_6_23_r2 = 1'b0;
logic din_almost_full_6_23;
assign din_6_23_r2.data   = 0;
assign din_6_23_r2.last   = 1'b0;
assign din_6_23_r2.bucket = 6;
rule_s_t din_6_24_r2;
logic din_valid_6_24_r2 = 1'b0;
logic din_almost_full_6_24;
assign din_6_24_r2.data   = 0;
assign din_6_24_r2.last   = 1'b0;
assign din_6_24_r2.bucket = 6;
rule_s_t din_6_25_r2;
logic din_valid_6_25_r2 = 1'b0;
logic din_almost_full_6_25;
assign din_6_25_r2.data   = 0;
assign din_6_25_r2.last   = 1'b0;
assign din_6_25_r2.bucket = 6;
rule_s_t din_6_26_r2;
logic din_valid_6_26_r2 = 1'b0;
logic din_almost_full_6_26;
assign din_6_26_r2.data   = 0;
assign din_6_26_r2.last   = 1'b0;
assign din_6_26_r2.bucket = 6;
rule_s_t din_6_27_r2;
logic din_valid_6_27_r2 = 1'b0;
logic din_almost_full_6_27;
assign din_6_27_r2.data   = 0;
assign din_6_27_r2.last   = 1'b0;
assign din_6_27_r2.bucket = 6;
rule_s_t din_6_28_r2;
logic din_valid_6_28_r2 = 1'b0;
logic din_almost_full_6_28;
assign din_6_28_r2.data   = 0;
assign din_6_28_r2.last   = 1'b0;
assign din_6_28_r2.bucket = 6;
rule_s_t din_6_29_r2;
logic din_valid_6_29_r2 = 1'b0;
logic din_almost_full_6_29;
assign din_6_29_r2.data   = 0;
assign din_6_29_r2.last   = 1'b0;
assign din_6_29_r2.bucket = 6;
rule_s_t din_6_30_r2;
logic din_valid_6_30_r2 = 1'b0;
logic din_almost_full_6_30;
assign din_6_30_r2.data   = 0;
assign din_6_30_r2.last   = 1'b0;
assign din_6_30_r2.bucket = 6;
rule_s_t din_6_31_r2;
logic din_valid_6_31_r2 = 1'b0;
logic din_almost_full_6_31;
assign din_6_31_r2.data   = 0;
assign din_6_31_r2.last   = 1'b0;
assign din_6_31_r2.bucket = 6;

logic [RID_WIDTH-1:0] hash_out_7_0;
logic hash_out_valid_filter_7_0;
rule_s_t din_7_0;
rule_s_t din_7_0_r1;
rule_s_t din_7_0_r2;
logic din_valid_7_0;
logic din_valid_7_0_r1;
logic din_valid_7_0_r2;
logic din_almost_full_7_0;
logic [RID_WIDTH-1:0] hash_out_7_1;
logic hash_out_valid_filter_7_1;
rule_s_t din_7_1;
rule_s_t din_7_1_r1;
rule_s_t din_7_1_r2;
logic din_valid_7_1;
logic din_valid_7_1_r1;
logic din_valid_7_1_r2;
logic din_almost_full_7_1;
logic [RID_WIDTH-1:0] hash_out_7_2;
logic hash_out_valid_filter_7_2;
rule_s_t din_7_2;
rule_s_t din_7_2_r1;
rule_s_t din_7_2_r2;
logic din_valid_7_2;
logic din_valid_7_2_r1;
logic din_valid_7_2_r2;
logic din_almost_full_7_2;
logic [RID_WIDTH-1:0] hash_out_7_3;
logic hash_out_valid_filter_7_3;
rule_s_t din_7_3;
rule_s_t din_7_3_r1;
rule_s_t din_7_3_r2;
logic din_valid_7_3;
logic din_valid_7_3_r1;
logic din_valid_7_3_r2;
logic din_almost_full_7_3;
logic [RID_WIDTH-1:0] hash_out_7_4;
logic hash_out_valid_filter_7_4;
rule_s_t din_7_4;
rule_s_t din_7_4_r1;
rule_s_t din_7_4_r2;
logic din_valid_7_4;
logic din_valid_7_4_r1;
logic din_valid_7_4_r2;
logic din_almost_full_7_4;
logic [RID_WIDTH-1:0] hash_out_7_5;
logic hash_out_valid_filter_7_5;
rule_s_t din_7_5;
rule_s_t din_7_5_r1;
rule_s_t din_7_5_r2;
logic din_valid_7_5;
logic din_valid_7_5_r1;
logic din_valid_7_5_r2;
logic din_almost_full_7_5;
logic [RID_WIDTH-1:0] hash_out_7_6;
logic hash_out_valid_filter_7_6;
rule_s_t din_7_6;
rule_s_t din_7_6_r1;
rule_s_t din_7_6_r2;
logic din_valid_7_6;
logic din_valid_7_6_r1;
logic din_valid_7_6_r2;
logic din_almost_full_7_6;
logic [RID_WIDTH-1:0] hash_out_7_7;
logic hash_out_valid_filter_7_7;
rule_s_t din_7_7;
rule_s_t din_7_7_r1;
rule_s_t din_7_7_r2;
logic din_valid_7_7;
logic din_valid_7_7_r1;
logic din_valid_7_7_r2;
logic din_almost_full_7_7;

rule_s_t din_7_8_r2;
logic din_valid_7_8_r2 = 1'b0;
logic din_almost_full_7_8;
assign din_7_8_r2.data   = 0;
assign din_7_8_r2.last   = 1'b0;
assign din_7_8_r2.bucket = 7;
rule_s_t din_7_9_r2;
logic din_valid_7_9_r2 = 1'b0;
logic din_almost_full_7_9;
assign din_7_9_r2.data   = 0;
assign din_7_9_r2.last   = 1'b0;
assign din_7_9_r2.bucket = 7;
rule_s_t din_7_10_r2;
logic din_valid_7_10_r2 = 1'b0;
logic din_almost_full_7_10;
assign din_7_10_r2.data   = 0;
assign din_7_10_r2.last   = 1'b0;
assign din_7_10_r2.bucket = 7;
rule_s_t din_7_11_r2;
logic din_valid_7_11_r2 = 1'b0;
logic din_almost_full_7_11;
assign din_7_11_r2.data   = 0;
assign din_7_11_r2.last   = 1'b0;
assign din_7_11_r2.bucket = 7;
rule_s_t din_7_12_r2;
logic din_valid_7_12_r2 = 1'b0;
logic din_almost_full_7_12;
assign din_7_12_r2.data   = 0;
assign din_7_12_r2.last   = 1'b0;
assign din_7_12_r2.bucket = 7;
rule_s_t din_7_13_r2;
logic din_valid_7_13_r2 = 1'b0;
logic din_almost_full_7_13;
assign din_7_13_r2.data   = 0;
assign din_7_13_r2.last   = 1'b0;
assign din_7_13_r2.bucket = 7;
rule_s_t din_7_14_r2;
logic din_valid_7_14_r2 = 1'b0;
logic din_almost_full_7_14;
assign din_7_14_r2.data   = 0;
assign din_7_14_r2.last   = 1'b0;
assign din_7_14_r2.bucket = 7;
rule_s_t din_7_15_r2;
logic din_valid_7_15_r2 = 1'b0;
logic din_almost_full_7_15;
assign din_7_15_r2.data   = 0;
assign din_7_15_r2.last   = 1'b0;
assign din_7_15_r2.bucket = 7;
rule_s_t din_7_16_r2;
logic din_valid_7_16_r2 = 1'b0;
logic din_almost_full_7_16;
assign din_7_16_r2.data   = 0;
assign din_7_16_r2.last   = 1'b0;
assign din_7_16_r2.bucket = 7;
rule_s_t din_7_17_r2;
logic din_valid_7_17_r2 = 1'b0;
logic din_almost_full_7_17;
assign din_7_17_r2.data   = 0;
assign din_7_17_r2.last   = 1'b0;
assign din_7_17_r2.bucket = 7;
rule_s_t din_7_18_r2;
logic din_valid_7_18_r2 = 1'b0;
logic din_almost_full_7_18;
assign din_7_18_r2.data   = 0;
assign din_7_18_r2.last   = 1'b0;
assign din_7_18_r2.bucket = 7;
rule_s_t din_7_19_r2;
logic din_valid_7_19_r2 = 1'b0;
logic din_almost_full_7_19;
assign din_7_19_r2.data   = 0;
assign din_7_19_r2.last   = 1'b0;
assign din_7_19_r2.bucket = 7;
rule_s_t din_7_20_r2;
logic din_valid_7_20_r2 = 1'b0;
logic din_almost_full_7_20;
assign din_7_20_r2.data   = 0;
assign din_7_20_r2.last   = 1'b0;
assign din_7_20_r2.bucket = 7;
rule_s_t din_7_21_r2;
logic din_valid_7_21_r2 = 1'b0;
logic din_almost_full_7_21;
assign din_7_21_r2.data   = 0;
assign din_7_21_r2.last   = 1'b0;
assign din_7_21_r2.bucket = 7;
rule_s_t din_7_22_r2;
logic din_valid_7_22_r2 = 1'b0;
logic din_almost_full_7_22;
assign din_7_22_r2.data   = 0;
assign din_7_22_r2.last   = 1'b0;
assign din_7_22_r2.bucket = 7;
rule_s_t din_7_23_r2;
logic din_valid_7_23_r2 = 1'b0;
logic din_almost_full_7_23;
assign din_7_23_r2.data   = 0;
assign din_7_23_r2.last   = 1'b0;
assign din_7_23_r2.bucket = 7;
rule_s_t din_7_24_r2;
logic din_valid_7_24_r2 = 1'b0;
logic din_almost_full_7_24;
assign din_7_24_r2.data   = 0;
assign din_7_24_r2.last   = 1'b0;
assign din_7_24_r2.bucket = 7;
rule_s_t din_7_25_r2;
logic din_valid_7_25_r2 = 1'b0;
logic din_almost_full_7_25;
assign din_7_25_r2.data   = 0;
assign din_7_25_r2.last   = 1'b0;
assign din_7_25_r2.bucket = 7;
rule_s_t din_7_26_r2;
logic din_valid_7_26_r2 = 1'b0;
logic din_almost_full_7_26;
assign din_7_26_r2.data   = 0;
assign din_7_26_r2.last   = 1'b0;
assign din_7_26_r2.bucket = 7;
rule_s_t din_7_27_r2;
logic din_valid_7_27_r2 = 1'b0;
logic din_almost_full_7_27;
assign din_7_27_r2.data   = 0;
assign din_7_27_r2.last   = 1'b0;
assign din_7_27_r2.bucket = 7;
rule_s_t din_7_28_r2;
logic din_valid_7_28_r2 = 1'b0;
logic din_almost_full_7_28;
assign din_7_28_r2.data   = 0;
assign din_7_28_r2.last   = 1'b0;
assign din_7_28_r2.bucket = 7;
rule_s_t din_7_29_r2;
logic din_valid_7_29_r2 = 1'b0;
logic din_almost_full_7_29;
assign din_7_29_r2.data   = 0;
assign din_7_29_r2.last   = 1'b0;
assign din_7_29_r2.bucket = 7;
rule_s_t din_7_30_r2;
logic din_valid_7_30_r2 = 1'b0;
logic din_almost_full_7_30;
assign din_7_30_r2.data   = 0;
assign din_7_30_r2.last   = 1'b0;
assign din_7_30_r2.bucket = 7;
rule_s_t din_7_31_r2;
logic din_valid_7_31_r2 = 1'b0;
logic din_almost_full_7_31;
assign din_7_31_r2.data   = 0;
assign din_7_31_r2.last   = 1'b0;
assign din_7_31_r2.bucket = 7;


logic out_new_pkt;

logic [255:0] in_convt;

assign in_convt[7+0*8:0+0*8] = in_data[255-0*8:255-7-0*8];
assign in_convt[7+1*8:0+1*8] = in_data[255-1*8:255-7-1*8];
assign in_convt[7+2*8:0+2*8] = in_data[255-2*8:255-7-2*8];
assign in_convt[7+3*8:0+3*8] = in_data[255-3*8:255-7-3*8];
assign in_convt[7+4*8:0+4*8] = in_data[255-4*8:255-7-4*8];
assign in_convt[7+5*8:0+5*8] = in_data[255-5*8:255-7-5*8];
assign in_convt[7+6*8:0+6*8] = in_data[255-6*8:255-7-6*8];
assign in_convt[7+7*8:0+7*8] = in_data[255-7*8:255-7-7*8];

always @ (posedge clk) begin
    in_ready <=   !din_almost_full_0_0 &  !din_almost_full_0_1 &  !din_almost_full_0_2 &  !din_almost_full_0_3 &  !din_almost_full_0_4 &  !din_almost_full_0_5 &  !din_almost_full_0_6 &  !din_almost_full_0_7 &    !din_almost_full_1_0 &  !din_almost_full_1_1 &  !din_almost_full_1_2 &  !din_almost_full_1_3 &  !din_almost_full_1_4 &  !din_almost_full_1_5 &  !din_almost_full_1_6 &  !din_almost_full_1_7 &    !din_almost_full_2_0 &  !din_almost_full_2_1 &  !din_almost_full_2_2 &  !din_almost_full_2_3 &  !din_almost_full_2_4 &  !din_almost_full_2_5 &  !din_almost_full_2_6 &  !din_almost_full_2_7 &    !din_almost_full_3_0 &  !din_almost_full_3_1 &  !din_almost_full_3_2 &  !din_almost_full_3_3 &  !din_almost_full_3_4 &  !din_almost_full_3_5 &  !din_almost_full_3_6 &  !din_almost_full_3_7 &    !din_almost_full_4_0 &  !din_almost_full_4_1 &  !din_almost_full_4_2 &  !din_almost_full_4_3 &  !din_almost_full_4_4 &  !din_almost_full_4_5 &  !din_almost_full_4_6 &  !din_almost_full_4_7 &    !din_almost_full_5_0 &  !din_almost_full_5_1 &  !din_almost_full_5_2 &  !din_almost_full_5_3 &  !din_almost_full_5_4 &  !din_almost_full_5_5 &  !din_almost_full_5_6 &  !din_almost_full_5_7 &    !din_almost_full_6_0 &  !din_almost_full_6_1 &  !din_almost_full_6_2 &  !din_almost_full_6_3 &  !din_almost_full_6_4 &  !din_almost_full_6_5 &  !din_almost_full_6_6 &  !din_almost_full_6_7 &    !din_almost_full_7_0 &  !din_almost_full_7_1 &  !din_almost_full_7_2 &  !din_almost_full_7_3 &  !din_almost_full_7_4 &  !din_almost_full_7_5 &  !din_almost_full_7_6 &  !din_almost_full_7_7 &   1;
    
    in_data_r1 <= in_convt;
    in_data_r2 <= in_data_r1;

    //only valid when the input is dequeued. 
    in_valid_r1 <= in_valid;
    in_valid_r2 <= in_valid_r1;
    init_r1 <= init;
    init_r2 <= init_r1;
    in_last_r1 <= in_last;
    in_last_r2 <= in_last_r1;
    in_strb_r1 <= in_strb;
    in_strb_r2 <= in_strb_r1;
end

always@(posedge clk)begin
    din_valid_0_0 <= out_new_pkt | hash_out_valid_filter_0_0;
    din_valid_0_0_r1 <= din_valid_0_0;
    din_valid_0_0_r2 <= din_valid_0_0_r1;

    din_0_0.data <= hash_out_valid_filter_0_0 ? hash_out_0_0 : 0;
    din_0_0.last <= out_new_pkt;
    din_0_0.bucket <= 0;


    din_0_0_r1 <= din_0_0;
    din_0_0_r2 <= din_0_0_r1;
    din_valid_0_1 <= out_new_pkt | hash_out_valid_filter_0_1;
    din_valid_0_1_r1 <= din_valid_0_1;
    din_valid_0_1_r2 <= din_valid_0_1_r1;

    din_0_1.data <= hash_out_valid_filter_0_1 ? hash_out_0_1 : 0;
    din_0_1.last <= out_new_pkt;
    din_0_1.bucket <= 0;


    din_0_1_r1 <= din_0_1;
    din_0_1_r2 <= din_0_1_r1;
    din_valid_0_2 <= out_new_pkt | hash_out_valid_filter_0_2;
    din_valid_0_2_r1 <= din_valid_0_2;
    din_valid_0_2_r2 <= din_valid_0_2_r1;

    din_0_2.data <= hash_out_valid_filter_0_2 ? hash_out_0_2 : 0;
    din_0_2.last <= out_new_pkt;
    din_0_2.bucket <= 0;


    din_0_2_r1 <= din_0_2;
    din_0_2_r2 <= din_0_2_r1;
    din_valid_0_3 <= out_new_pkt | hash_out_valid_filter_0_3;
    din_valid_0_3_r1 <= din_valid_0_3;
    din_valid_0_3_r2 <= din_valid_0_3_r1;

    din_0_3.data <= hash_out_valid_filter_0_3 ? hash_out_0_3 : 0;
    din_0_3.last <= out_new_pkt;
    din_0_3.bucket <= 0;


    din_0_3_r1 <= din_0_3;
    din_0_3_r2 <= din_0_3_r1;
    din_valid_0_4 <= out_new_pkt | hash_out_valid_filter_0_4;
    din_valid_0_4_r1 <= din_valid_0_4;
    din_valid_0_4_r2 <= din_valid_0_4_r1;

    din_0_4.data <= hash_out_valid_filter_0_4 ? hash_out_0_4 : 0;
    din_0_4.last <= out_new_pkt;
    din_0_4.bucket <= 0;


    din_0_4_r1 <= din_0_4;
    din_0_4_r2 <= din_0_4_r1;
    din_valid_0_5 <= out_new_pkt | hash_out_valid_filter_0_5;
    din_valid_0_5_r1 <= din_valid_0_5;
    din_valid_0_5_r2 <= din_valid_0_5_r1;

    din_0_5.data <= hash_out_valid_filter_0_5 ? hash_out_0_5 : 0;
    din_0_5.last <= out_new_pkt;
    din_0_5.bucket <= 0;


    din_0_5_r1 <= din_0_5;
    din_0_5_r2 <= din_0_5_r1;
    din_valid_0_6 <= out_new_pkt | hash_out_valid_filter_0_6;
    din_valid_0_6_r1 <= din_valid_0_6;
    din_valid_0_6_r2 <= din_valid_0_6_r1;

    din_0_6.data <= hash_out_valid_filter_0_6 ? hash_out_0_6 : 0;
    din_0_6.last <= out_new_pkt;
    din_0_6.bucket <= 0;


    din_0_6_r1 <= din_0_6;
    din_0_6_r2 <= din_0_6_r1;
    din_valid_0_7 <= out_new_pkt | hash_out_valid_filter_0_7;
    din_valid_0_7_r1 <= din_valid_0_7;
    din_valid_0_7_r2 <= din_valid_0_7_r1;

    din_0_7.data <= hash_out_valid_filter_0_7 ? hash_out_0_7 : 0;
    din_0_7.last <= out_new_pkt;
    din_0_7.bucket <= 0;


    din_0_7_r1 <= din_0_7;
    din_0_7_r2 <= din_0_7_r1;
    din_valid_1_0 <= out_new_pkt | hash_out_valid_filter_1_0;
    din_valid_1_0_r1 <= din_valid_1_0;
    din_valid_1_0_r2 <= din_valid_1_0_r1;

    din_1_0.data <= hash_out_valid_filter_1_0 ? hash_out_1_0 : 0;
    din_1_0.last <= out_new_pkt;
    din_1_0.bucket <= 1;


    din_1_0_r1 <= din_1_0;
    din_1_0_r2 <= din_1_0_r1;
    din_valid_1_1 <= out_new_pkt | hash_out_valid_filter_1_1;
    din_valid_1_1_r1 <= din_valid_1_1;
    din_valid_1_1_r2 <= din_valid_1_1_r1;

    din_1_1.data <= hash_out_valid_filter_1_1 ? hash_out_1_1 : 0;
    din_1_1.last <= out_new_pkt;
    din_1_1.bucket <= 1;


    din_1_1_r1 <= din_1_1;
    din_1_1_r2 <= din_1_1_r1;
    din_valid_1_2 <= out_new_pkt | hash_out_valid_filter_1_2;
    din_valid_1_2_r1 <= din_valid_1_2;
    din_valid_1_2_r2 <= din_valid_1_2_r1;

    din_1_2.data <= hash_out_valid_filter_1_2 ? hash_out_1_2 : 0;
    din_1_2.last <= out_new_pkt;
    din_1_2.bucket <= 1;


    din_1_2_r1 <= din_1_2;
    din_1_2_r2 <= din_1_2_r1;
    din_valid_1_3 <= out_new_pkt | hash_out_valid_filter_1_3;
    din_valid_1_3_r1 <= din_valid_1_3;
    din_valid_1_3_r2 <= din_valid_1_3_r1;

    din_1_3.data <= hash_out_valid_filter_1_3 ? hash_out_1_3 : 0;
    din_1_3.last <= out_new_pkt;
    din_1_3.bucket <= 1;


    din_1_3_r1 <= din_1_3;
    din_1_3_r2 <= din_1_3_r1;
    din_valid_1_4 <= out_new_pkt | hash_out_valid_filter_1_4;
    din_valid_1_4_r1 <= din_valid_1_4;
    din_valid_1_4_r2 <= din_valid_1_4_r1;

    din_1_4.data <= hash_out_valid_filter_1_4 ? hash_out_1_4 : 0;
    din_1_4.last <= out_new_pkt;
    din_1_4.bucket <= 1;


    din_1_4_r1 <= din_1_4;
    din_1_4_r2 <= din_1_4_r1;
    din_valid_1_5 <= out_new_pkt | hash_out_valid_filter_1_5;
    din_valid_1_5_r1 <= din_valid_1_5;
    din_valid_1_5_r2 <= din_valid_1_5_r1;

    din_1_5.data <= hash_out_valid_filter_1_5 ? hash_out_1_5 : 0;
    din_1_5.last <= out_new_pkt;
    din_1_5.bucket <= 1;


    din_1_5_r1 <= din_1_5;
    din_1_5_r2 <= din_1_5_r1;
    din_valid_1_6 <= out_new_pkt | hash_out_valid_filter_1_6;
    din_valid_1_6_r1 <= din_valid_1_6;
    din_valid_1_6_r2 <= din_valid_1_6_r1;

    din_1_6.data <= hash_out_valid_filter_1_6 ? hash_out_1_6 : 0;
    din_1_6.last <= out_new_pkt;
    din_1_6.bucket <= 1;


    din_1_6_r1 <= din_1_6;
    din_1_6_r2 <= din_1_6_r1;
    din_valid_1_7 <= out_new_pkt | hash_out_valid_filter_1_7;
    din_valid_1_7_r1 <= din_valid_1_7;
    din_valid_1_7_r2 <= din_valid_1_7_r1;

    din_1_7.data <= hash_out_valid_filter_1_7 ? hash_out_1_7 : 0;
    din_1_7.last <= out_new_pkt;
    din_1_7.bucket <= 1;


    din_1_7_r1 <= din_1_7;
    din_1_7_r2 <= din_1_7_r1;
    din_valid_2_0 <= out_new_pkt | hash_out_valid_filter_2_0;
    din_valid_2_0_r1 <= din_valid_2_0;
    din_valid_2_0_r2 <= din_valid_2_0_r1;

    din_2_0.data <= hash_out_valid_filter_2_0 ? hash_out_2_0 : 0;
    din_2_0.last <= out_new_pkt;
    din_2_0.bucket <= 2;


    din_2_0_r1 <= din_2_0;
    din_2_0_r2 <= din_2_0_r1;
    din_valid_2_1 <= out_new_pkt | hash_out_valid_filter_2_1;
    din_valid_2_1_r1 <= din_valid_2_1;
    din_valid_2_1_r2 <= din_valid_2_1_r1;

    din_2_1.data <= hash_out_valid_filter_2_1 ? hash_out_2_1 : 0;
    din_2_1.last <= out_new_pkt;
    din_2_1.bucket <= 2;


    din_2_1_r1 <= din_2_1;
    din_2_1_r2 <= din_2_1_r1;
    din_valid_2_2 <= out_new_pkt | hash_out_valid_filter_2_2;
    din_valid_2_2_r1 <= din_valid_2_2;
    din_valid_2_2_r2 <= din_valid_2_2_r1;

    din_2_2.data <= hash_out_valid_filter_2_2 ? hash_out_2_2 : 0;
    din_2_2.last <= out_new_pkt;
    din_2_2.bucket <= 2;


    din_2_2_r1 <= din_2_2;
    din_2_2_r2 <= din_2_2_r1;
    din_valid_2_3 <= out_new_pkt | hash_out_valid_filter_2_3;
    din_valid_2_3_r1 <= din_valid_2_3;
    din_valid_2_3_r2 <= din_valid_2_3_r1;

    din_2_3.data <= hash_out_valid_filter_2_3 ? hash_out_2_3 : 0;
    din_2_3.last <= out_new_pkt;
    din_2_3.bucket <= 2;


    din_2_3_r1 <= din_2_3;
    din_2_3_r2 <= din_2_3_r1;
    din_valid_2_4 <= out_new_pkt | hash_out_valid_filter_2_4;
    din_valid_2_4_r1 <= din_valid_2_4;
    din_valid_2_4_r2 <= din_valid_2_4_r1;

    din_2_4.data <= hash_out_valid_filter_2_4 ? hash_out_2_4 : 0;
    din_2_4.last <= out_new_pkt;
    din_2_4.bucket <= 2;


    din_2_4_r1 <= din_2_4;
    din_2_4_r2 <= din_2_4_r1;
    din_valid_2_5 <= out_new_pkt | hash_out_valid_filter_2_5;
    din_valid_2_5_r1 <= din_valid_2_5;
    din_valid_2_5_r2 <= din_valid_2_5_r1;

    din_2_5.data <= hash_out_valid_filter_2_5 ? hash_out_2_5 : 0;
    din_2_5.last <= out_new_pkt;
    din_2_5.bucket <= 2;


    din_2_5_r1 <= din_2_5;
    din_2_5_r2 <= din_2_5_r1;
    din_valid_2_6 <= out_new_pkt | hash_out_valid_filter_2_6;
    din_valid_2_6_r1 <= din_valid_2_6;
    din_valid_2_6_r2 <= din_valid_2_6_r1;

    din_2_6.data <= hash_out_valid_filter_2_6 ? hash_out_2_6 : 0;
    din_2_6.last <= out_new_pkt;
    din_2_6.bucket <= 2;


    din_2_6_r1 <= din_2_6;
    din_2_6_r2 <= din_2_6_r1;
    din_valid_2_7 <= out_new_pkt | hash_out_valid_filter_2_7;
    din_valid_2_7_r1 <= din_valid_2_7;
    din_valid_2_7_r2 <= din_valid_2_7_r1;

    din_2_7.data <= hash_out_valid_filter_2_7 ? hash_out_2_7 : 0;
    din_2_7.last <= out_new_pkt;
    din_2_7.bucket <= 2;


    din_2_7_r1 <= din_2_7;
    din_2_7_r2 <= din_2_7_r1;
    din_valid_3_0 <= out_new_pkt | hash_out_valid_filter_3_0;
    din_valid_3_0_r1 <= din_valid_3_0;
    din_valid_3_0_r2 <= din_valid_3_0_r1;

    din_3_0.data <= hash_out_valid_filter_3_0 ? hash_out_3_0 : 0;
    din_3_0.last <= out_new_pkt;
    din_3_0.bucket <= 3;


    din_3_0_r1 <= din_3_0;
    din_3_0_r2 <= din_3_0_r1;
    din_valid_3_1 <= out_new_pkt | hash_out_valid_filter_3_1;
    din_valid_3_1_r1 <= din_valid_3_1;
    din_valid_3_1_r2 <= din_valid_3_1_r1;

    din_3_1.data <= hash_out_valid_filter_3_1 ? hash_out_3_1 : 0;
    din_3_1.last <= out_new_pkt;
    din_3_1.bucket <= 3;


    din_3_1_r1 <= din_3_1;
    din_3_1_r2 <= din_3_1_r1;
    din_valid_3_2 <= out_new_pkt | hash_out_valid_filter_3_2;
    din_valid_3_2_r1 <= din_valid_3_2;
    din_valid_3_2_r2 <= din_valid_3_2_r1;

    din_3_2.data <= hash_out_valid_filter_3_2 ? hash_out_3_2 : 0;
    din_3_2.last <= out_new_pkt;
    din_3_2.bucket <= 3;


    din_3_2_r1 <= din_3_2;
    din_3_2_r2 <= din_3_2_r1;
    din_valid_3_3 <= out_new_pkt | hash_out_valid_filter_3_3;
    din_valid_3_3_r1 <= din_valid_3_3;
    din_valid_3_3_r2 <= din_valid_3_3_r1;

    din_3_3.data <= hash_out_valid_filter_3_3 ? hash_out_3_3 : 0;
    din_3_3.last <= out_new_pkt;
    din_3_3.bucket <= 3;


    din_3_3_r1 <= din_3_3;
    din_3_3_r2 <= din_3_3_r1;
    din_valid_3_4 <= out_new_pkt | hash_out_valid_filter_3_4;
    din_valid_3_4_r1 <= din_valid_3_4;
    din_valid_3_4_r2 <= din_valid_3_4_r1;

    din_3_4.data <= hash_out_valid_filter_3_4 ? hash_out_3_4 : 0;
    din_3_4.last <= out_new_pkt;
    din_3_4.bucket <= 3;


    din_3_4_r1 <= din_3_4;
    din_3_4_r2 <= din_3_4_r1;
    din_valid_3_5 <= out_new_pkt | hash_out_valid_filter_3_5;
    din_valid_3_5_r1 <= din_valid_3_5;
    din_valid_3_5_r2 <= din_valid_3_5_r1;

    din_3_5.data <= hash_out_valid_filter_3_5 ? hash_out_3_5 : 0;
    din_3_5.last <= out_new_pkt;
    din_3_5.bucket <= 3;


    din_3_5_r1 <= din_3_5;
    din_3_5_r2 <= din_3_5_r1;
    din_valid_3_6 <= out_new_pkt | hash_out_valid_filter_3_6;
    din_valid_3_6_r1 <= din_valid_3_6;
    din_valid_3_6_r2 <= din_valid_3_6_r1;

    din_3_6.data <= hash_out_valid_filter_3_6 ? hash_out_3_6 : 0;
    din_3_6.last <= out_new_pkt;
    din_3_6.bucket <= 3;


    din_3_6_r1 <= din_3_6;
    din_3_6_r2 <= din_3_6_r1;
    din_valid_3_7 <= out_new_pkt | hash_out_valid_filter_3_7;
    din_valid_3_7_r1 <= din_valid_3_7;
    din_valid_3_7_r2 <= din_valid_3_7_r1;

    din_3_7.data <= hash_out_valid_filter_3_7 ? hash_out_3_7 : 0;
    din_3_7.last <= out_new_pkt;
    din_3_7.bucket <= 3;


    din_3_7_r1 <= din_3_7;
    din_3_7_r2 <= din_3_7_r1;
    din_valid_4_0 <= out_new_pkt | hash_out_valid_filter_4_0;
    din_valid_4_0_r1 <= din_valid_4_0;
    din_valid_4_0_r2 <= din_valid_4_0_r1;

    din_4_0.data <= hash_out_valid_filter_4_0 ? hash_out_4_0 : 0;
    din_4_0.last <= out_new_pkt;
    din_4_0.bucket <= 4;


    din_4_0_r1 <= din_4_0;
    din_4_0_r2 <= din_4_0_r1;
    din_valid_4_1 <= out_new_pkt | hash_out_valid_filter_4_1;
    din_valid_4_1_r1 <= din_valid_4_1;
    din_valid_4_1_r2 <= din_valid_4_1_r1;

    din_4_1.data <= hash_out_valid_filter_4_1 ? hash_out_4_1 : 0;
    din_4_1.last <= out_new_pkt;
    din_4_1.bucket <= 4;


    din_4_1_r1 <= din_4_1;
    din_4_1_r2 <= din_4_1_r1;
    din_valid_4_2 <= out_new_pkt | hash_out_valid_filter_4_2;
    din_valid_4_2_r1 <= din_valid_4_2;
    din_valid_4_2_r2 <= din_valid_4_2_r1;

    din_4_2.data <= hash_out_valid_filter_4_2 ? hash_out_4_2 : 0;
    din_4_2.last <= out_new_pkt;
    din_4_2.bucket <= 4;


    din_4_2_r1 <= din_4_2;
    din_4_2_r2 <= din_4_2_r1;
    din_valid_4_3 <= out_new_pkt | hash_out_valid_filter_4_3;
    din_valid_4_3_r1 <= din_valid_4_3;
    din_valid_4_3_r2 <= din_valid_4_3_r1;

    din_4_3.data <= hash_out_valid_filter_4_3 ? hash_out_4_3 : 0;
    din_4_3.last <= out_new_pkt;
    din_4_3.bucket <= 4;


    din_4_3_r1 <= din_4_3;
    din_4_3_r2 <= din_4_3_r1;
    din_valid_4_4 <= out_new_pkt | hash_out_valid_filter_4_4;
    din_valid_4_4_r1 <= din_valid_4_4;
    din_valid_4_4_r2 <= din_valid_4_4_r1;

    din_4_4.data <= hash_out_valid_filter_4_4 ? hash_out_4_4 : 0;
    din_4_4.last <= out_new_pkt;
    din_4_4.bucket <= 4;


    din_4_4_r1 <= din_4_4;
    din_4_4_r2 <= din_4_4_r1;
    din_valid_4_5 <= out_new_pkt | hash_out_valid_filter_4_5;
    din_valid_4_5_r1 <= din_valid_4_5;
    din_valid_4_5_r2 <= din_valid_4_5_r1;

    din_4_5.data <= hash_out_valid_filter_4_5 ? hash_out_4_5 : 0;
    din_4_5.last <= out_new_pkt;
    din_4_5.bucket <= 4;


    din_4_5_r1 <= din_4_5;
    din_4_5_r2 <= din_4_5_r1;
    din_valid_4_6 <= out_new_pkt | hash_out_valid_filter_4_6;
    din_valid_4_6_r1 <= din_valid_4_6;
    din_valid_4_6_r2 <= din_valid_4_6_r1;

    din_4_6.data <= hash_out_valid_filter_4_6 ? hash_out_4_6 : 0;
    din_4_6.last <= out_new_pkt;
    din_4_6.bucket <= 4;


    din_4_6_r1 <= din_4_6;
    din_4_6_r2 <= din_4_6_r1;
    din_valid_4_7 <= out_new_pkt | hash_out_valid_filter_4_7;
    din_valid_4_7_r1 <= din_valid_4_7;
    din_valid_4_7_r2 <= din_valid_4_7_r1;

    din_4_7.data <= hash_out_valid_filter_4_7 ? hash_out_4_7 : 0;
    din_4_7.last <= out_new_pkt;
    din_4_7.bucket <= 4;


    din_4_7_r1 <= din_4_7;
    din_4_7_r2 <= din_4_7_r1;
    din_valid_5_0 <= out_new_pkt | hash_out_valid_filter_5_0;
    din_valid_5_0_r1 <= din_valid_5_0;
    din_valid_5_0_r2 <= din_valid_5_0_r1;

    din_5_0.data <= hash_out_valid_filter_5_0 ? hash_out_5_0 : 0;
    din_5_0.last <= out_new_pkt;
    din_5_0.bucket <= 5;


    din_5_0_r1 <= din_5_0;
    din_5_0_r2 <= din_5_0_r1;
    din_valid_5_1 <= out_new_pkt | hash_out_valid_filter_5_1;
    din_valid_5_1_r1 <= din_valid_5_1;
    din_valid_5_1_r2 <= din_valid_5_1_r1;

    din_5_1.data <= hash_out_valid_filter_5_1 ? hash_out_5_1 : 0;
    din_5_1.last <= out_new_pkt;
    din_5_1.bucket <= 5;


    din_5_1_r1 <= din_5_1;
    din_5_1_r2 <= din_5_1_r1;
    din_valid_5_2 <= out_new_pkt | hash_out_valid_filter_5_2;
    din_valid_5_2_r1 <= din_valid_5_2;
    din_valid_5_2_r2 <= din_valid_5_2_r1;

    din_5_2.data <= hash_out_valid_filter_5_2 ? hash_out_5_2 : 0;
    din_5_2.last <= out_new_pkt;
    din_5_2.bucket <= 5;


    din_5_2_r1 <= din_5_2;
    din_5_2_r2 <= din_5_2_r1;
    din_valid_5_3 <= out_new_pkt | hash_out_valid_filter_5_3;
    din_valid_5_3_r1 <= din_valid_5_3;
    din_valid_5_3_r2 <= din_valid_5_3_r1;

    din_5_3.data <= hash_out_valid_filter_5_3 ? hash_out_5_3 : 0;
    din_5_3.last <= out_new_pkt;
    din_5_3.bucket <= 5;


    din_5_3_r1 <= din_5_3;
    din_5_3_r2 <= din_5_3_r1;
    din_valid_5_4 <= out_new_pkt | hash_out_valid_filter_5_4;
    din_valid_5_4_r1 <= din_valid_5_4;
    din_valid_5_4_r2 <= din_valid_5_4_r1;

    din_5_4.data <= hash_out_valid_filter_5_4 ? hash_out_5_4 : 0;
    din_5_4.last <= out_new_pkt;
    din_5_4.bucket <= 5;


    din_5_4_r1 <= din_5_4;
    din_5_4_r2 <= din_5_4_r1;
    din_valid_5_5 <= out_new_pkt | hash_out_valid_filter_5_5;
    din_valid_5_5_r1 <= din_valid_5_5;
    din_valid_5_5_r2 <= din_valid_5_5_r1;

    din_5_5.data <= hash_out_valid_filter_5_5 ? hash_out_5_5 : 0;
    din_5_5.last <= out_new_pkt;
    din_5_5.bucket <= 5;


    din_5_5_r1 <= din_5_5;
    din_5_5_r2 <= din_5_5_r1;
    din_valid_5_6 <= out_new_pkt | hash_out_valid_filter_5_6;
    din_valid_5_6_r1 <= din_valid_5_6;
    din_valid_5_6_r2 <= din_valid_5_6_r1;

    din_5_6.data <= hash_out_valid_filter_5_6 ? hash_out_5_6 : 0;
    din_5_6.last <= out_new_pkt;
    din_5_6.bucket <= 5;


    din_5_6_r1 <= din_5_6;
    din_5_6_r2 <= din_5_6_r1;
    din_valid_5_7 <= out_new_pkt | hash_out_valid_filter_5_7;
    din_valid_5_7_r1 <= din_valid_5_7;
    din_valid_5_7_r2 <= din_valid_5_7_r1;

    din_5_7.data <= hash_out_valid_filter_5_7 ? hash_out_5_7 : 0;
    din_5_7.last <= out_new_pkt;
    din_5_7.bucket <= 5;


    din_5_7_r1 <= din_5_7;
    din_5_7_r2 <= din_5_7_r1;
    din_valid_6_0 <= out_new_pkt | hash_out_valid_filter_6_0;
    din_valid_6_0_r1 <= din_valid_6_0;
    din_valid_6_0_r2 <= din_valid_6_0_r1;

    din_6_0.data <= hash_out_valid_filter_6_0 ? hash_out_6_0 : 0;
    din_6_0.last <= out_new_pkt;
    din_6_0.bucket <= 6;


    din_6_0_r1 <= din_6_0;
    din_6_0_r2 <= din_6_0_r1;
    din_valid_6_1 <= out_new_pkt | hash_out_valid_filter_6_1;
    din_valid_6_1_r1 <= din_valid_6_1;
    din_valid_6_1_r2 <= din_valid_6_1_r1;

    din_6_1.data <= hash_out_valid_filter_6_1 ? hash_out_6_1 : 0;
    din_6_1.last <= out_new_pkt;
    din_6_1.bucket <= 6;


    din_6_1_r1 <= din_6_1;
    din_6_1_r2 <= din_6_1_r1;
    din_valid_6_2 <= out_new_pkt | hash_out_valid_filter_6_2;
    din_valid_6_2_r1 <= din_valid_6_2;
    din_valid_6_2_r2 <= din_valid_6_2_r1;

    din_6_2.data <= hash_out_valid_filter_6_2 ? hash_out_6_2 : 0;
    din_6_2.last <= out_new_pkt;
    din_6_2.bucket <= 6;


    din_6_2_r1 <= din_6_2;
    din_6_2_r2 <= din_6_2_r1;
    din_valid_6_3 <= out_new_pkt | hash_out_valid_filter_6_3;
    din_valid_6_3_r1 <= din_valid_6_3;
    din_valid_6_3_r2 <= din_valid_6_3_r1;

    din_6_3.data <= hash_out_valid_filter_6_3 ? hash_out_6_3 : 0;
    din_6_3.last <= out_new_pkt;
    din_6_3.bucket <= 6;


    din_6_3_r1 <= din_6_3;
    din_6_3_r2 <= din_6_3_r1;
    din_valid_6_4 <= out_new_pkt | hash_out_valid_filter_6_4;
    din_valid_6_4_r1 <= din_valid_6_4;
    din_valid_6_4_r2 <= din_valid_6_4_r1;

    din_6_4.data <= hash_out_valid_filter_6_4 ? hash_out_6_4 : 0;
    din_6_4.last <= out_new_pkt;
    din_6_4.bucket <= 6;


    din_6_4_r1 <= din_6_4;
    din_6_4_r2 <= din_6_4_r1;
    din_valid_6_5 <= out_new_pkt | hash_out_valid_filter_6_5;
    din_valid_6_5_r1 <= din_valid_6_5;
    din_valid_6_5_r2 <= din_valid_6_5_r1;

    din_6_5.data <= hash_out_valid_filter_6_5 ? hash_out_6_5 : 0;
    din_6_5.last <= out_new_pkt;
    din_6_5.bucket <= 6;


    din_6_5_r1 <= din_6_5;
    din_6_5_r2 <= din_6_5_r1;
    din_valid_6_6 <= out_new_pkt | hash_out_valid_filter_6_6;
    din_valid_6_6_r1 <= din_valid_6_6;
    din_valid_6_6_r2 <= din_valid_6_6_r1;

    din_6_6.data <= hash_out_valid_filter_6_6 ? hash_out_6_6 : 0;
    din_6_6.last <= out_new_pkt;
    din_6_6.bucket <= 6;


    din_6_6_r1 <= din_6_6;
    din_6_6_r2 <= din_6_6_r1;
    din_valid_6_7 <= out_new_pkt | hash_out_valid_filter_6_7;
    din_valid_6_7_r1 <= din_valid_6_7;
    din_valid_6_7_r2 <= din_valid_6_7_r1;

    din_6_7.data <= hash_out_valid_filter_6_7 ? hash_out_6_7 : 0;
    din_6_7.last <= out_new_pkt;
    din_6_7.bucket <= 6;


    din_6_7_r1 <= din_6_7;
    din_6_7_r2 <= din_6_7_r1;
    din_valid_7_0 <= out_new_pkt | hash_out_valid_filter_7_0;
    din_valid_7_0_r1 <= din_valid_7_0;
    din_valid_7_0_r2 <= din_valid_7_0_r1;

    din_7_0.data <= hash_out_valid_filter_7_0 ? hash_out_7_0 : 0;
    din_7_0.last <= out_new_pkt;
    din_7_0.bucket <= 7;


    din_7_0_r1 <= din_7_0;
    din_7_0_r2 <= din_7_0_r1;
    din_valid_7_1 <= out_new_pkt | hash_out_valid_filter_7_1;
    din_valid_7_1_r1 <= din_valid_7_1;
    din_valid_7_1_r2 <= din_valid_7_1_r1;

    din_7_1.data <= hash_out_valid_filter_7_1 ? hash_out_7_1 : 0;
    din_7_1.last <= out_new_pkt;
    din_7_1.bucket <= 7;


    din_7_1_r1 <= din_7_1;
    din_7_1_r2 <= din_7_1_r1;
    din_valid_7_2 <= out_new_pkt | hash_out_valid_filter_7_2;
    din_valid_7_2_r1 <= din_valid_7_2;
    din_valid_7_2_r2 <= din_valid_7_2_r1;

    din_7_2.data <= hash_out_valid_filter_7_2 ? hash_out_7_2 : 0;
    din_7_2.last <= out_new_pkt;
    din_7_2.bucket <= 7;


    din_7_2_r1 <= din_7_2;
    din_7_2_r2 <= din_7_2_r1;
    din_valid_7_3 <= out_new_pkt | hash_out_valid_filter_7_3;
    din_valid_7_3_r1 <= din_valid_7_3;
    din_valid_7_3_r2 <= din_valid_7_3_r1;

    din_7_3.data <= hash_out_valid_filter_7_3 ? hash_out_7_3 : 0;
    din_7_3.last <= out_new_pkt;
    din_7_3.bucket <= 7;


    din_7_3_r1 <= din_7_3;
    din_7_3_r2 <= din_7_3_r1;
    din_valid_7_4 <= out_new_pkt | hash_out_valid_filter_7_4;
    din_valid_7_4_r1 <= din_valid_7_4;
    din_valid_7_4_r2 <= din_valid_7_4_r1;

    din_7_4.data <= hash_out_valid_filter_7_4 ? hash_out_7_4 : 0;
    din_7_4.last <= out_new_pkt;
    din_7_4.bucket <= 7;


    din_7_4_r1 <= din_7_4;
    din_7_4_r2 <= din_7_4_r1;
    din_valid_7_5 <= out_new_pkt | hash_out_valid_filter_7_5;
    din_valid_7_5_r1 <= din_valid_7_5;
    din_valid_7_5_r2 <= din_valid_7_5_r1;

    din_7_5.data <= hash_out_valid_filter_7_5 ? hash_out_7_5 : 0;
    din_7_5.last <= out_new_pkt;
    din_7_5.bucket <= 7;


    din_7_5_r1 <= din_7_5;
    din_7_5_r2 <= din_7_5_r1;
    din_valid_7_6 <= out_new_pkt | hash_out_valid_filter_7_6;
    din_valid_7_6_r1 <= din_valid_7_6;
    din_valid_7_6_r2 <= din_valid_7_6_r1;

    din_7_6.data <= hash_out_valid_filter_7_6 ? hash_out_7_6 : 0;
    din_7_6.last <= out_new_pkt;
    din_7_6.bucket <= 7;


    din_7_6_r1 <= din_7_6;
    din_7_6_r2 <= din_7_6_r1;
    din_valid_7_7 <= out_new_pkt | hash_out_valid_filter_7_7;
    din_valid_7_7_r1 <= din_valid_7_7;
    din_valid_7_7_r2 <= din_valid_7_7_r1;

    din_7_7.data <= hash_out_valid_filter_7_7 ? hash_out_7_7 : 0;
    din_7_7.last <= out_new_pkt;
    din_7_7.bucket <= 7;


    din_7_7_r1 <= din_7_7;
    din_7_7_r2 <= din_7_7_r1;
end

//Instantiation
frontend front(
    .clk(clk),
    .rst(rst),
    .hash_out_0_0(hash_out_0_0),
    .hash_out_valid_filter_0_0(hash_out_valid_filter_0_0),
    .hash_out_0_1(hash_out_0_1),
    .hash_out_valid_filter_0_1(hash_out_valid_filter_0_1),
    .hash_out_0_2(hash_out_0_2),
    .hash_out_valid_filter_0_2(hash_out_valid_filter_0_2),
    .hash_out_0_3(hash_out_0_3),
    .hash_out_valid_filter_0_3(hash_out_valid_filter_0_3),
    .hash_out_0_4(hash_out_0_4),
    .hash_out_valid_filter_0_4(hash_out_valid_filter_0_4),
    .hash_out_0_5(hash_out_0_5),
    .hash_out_valid_filter_0_5(hash_out_valid_filter_0_5),
    .hash_out_0_6(hash_out_0_6),
    .hash_out_valid_filter_0_6(hash_out_valid_filter_0_6),
    .hash_out_0_7(hash_out_0_7),
    .hash_out_valid_filter_0_7(hash_out_valid_filter_0_7),
    .hash_out_1_0(hash_out_1_0),
    .hash_out_valid_filter_1_0(hash_out_valid_filter_1_0),
    .hash_out_1_1(hash_out_1_1),
    .hash_out_valid_filter_1_1(hash_out_valid_filter_1_1),
    .hash_out_1_2(hash_out_1_2),
    .hash_out_valid_filter_1_2(hash_out_valid_filter_1_2),
    .hash_out_1_3(hash_out_1_3),
    .hash_out_valid_filter_1_3(hash_out_valid_filter_1_3),
    .hash_out_1_4(hash_out_1_4),
    .hash_out_valid_filter_1_4(hash_out_valid_filter_1_4),
    .hash_out_1_5(hash_out_1_5),
    .hash_out_valid_filter_1_5(hash_out_valid_filter_1_5),
    .hash_out_1_6(hash_out_1_6),
    .hash_out_valid_filter_1_6(hash_out_valid_filter_1_6),
    .hash_out_1_7(hash_out_1_7),
    .hash_out_valid_filter_1_7(hash_out_valid_filter_1_7),
    .hash_out_2_0(hash_out_2_0),
    .hash_out_valid_filter_2_0(hash_out_valid_filter_2_0),
    .hash_out_2_1(hash_out_2_1),
    .hash_out_valid_filter_2_1(hash_out_valid_filter_2_1),
    .hash_out_2_2(hash_out_2_2),
    .hash_out_valid_filter_2_2(hash_out_valid_filter_2_2),
    .hash_out_2_3(hash_out_2_3),
    .hash_out_valid_filter_2_3(hash_out_valid_filter_2_3),
    .hash_out_2_4(hash_out_2_4),
    .hash_out_valid_filter_2_4(hash_out_valid_filter_2_4),
    .hash_out_2_5(hash_out_2_5),
    .hash_out_valid_filter_2_5(hash_out_valid_filter_2_5),
    .hash_out_2_6(hash_out_2_6),
    .hash_out_valid_filter_2_6(hash_out_valid_filter_2_6),
    .hash_out_2_7(hash_out_2_7),
    .hash_out_valid_filter_2_7(hash_out_valid_filter_2_7),
    .hash_out_3_0(hash_out_3_0),
    .hash_out_valid_filter_3_0(hash_out_valid_filter_3_0),
    .hash_out_3_1(hash_out_3_1),
    .hash_out_valid_filter_3_1(hash_out_valid_filter_3_1),
    .hash_out_3_2(hash_out_3_2),
    .hash_out_valid_filter_3_2(hash_out_valid_filter_3_2),
    .hash_out_3_3(hash_out_3_3),
    .hash_out_valid_filter_3_3(hash_out_valid_filter_3_3),
    .hash_out_3_4(hash_out_3_4),
    .hash_out_valid_filter_3_4(hash_out_valid_filter_3_4),
    .hash_out_3_5(hash_out_3_5),
    .hash_out_valid_filter_3_5(hash_out_valid_filter_3_5),
    .hash_out_3_6(hash_out_3_6),
    .hash_out_valid_filter_3_6(hash_out_valid_filter_3_6),
    .hash_out_3_7(hash_out_3_7),
    .hash_out_valid_filter_3_7(hash_out_valid_filter_3_7),
    .hash_out_4_0(hash_out_4_0),
    .hash_out_valid_filter_4_0(hash_out_valid_filter_4_0),
    .hash_out_4_1(hash_out_4_1),
    .hash_out_valid_filter_4_1(hash_out_valid_filter_4_1),
    .hash_out_4_2(hash_out_4_2),
    .hash_out_valid_filter_4_2(hash_out_valid_filter_4_2),
    .hash_out_4_3(hash_out_4_3),
    .hash_out_valid_filter_4_3(hash_out_valid_filter_4_3),
    .hash_out_4_4(hash_out_4_4),
    .hash_out_valid_filter_4_4(hash_out_valid_filter_4_4),
    .hash_out_4_5(hash_out_4_5),
    .hash_out_valid_filter_4_5(hash_out_valid_filter_4_5),
    .hash_out_4_6(hash_out_4_6),
    .hash_out_valid_filter_4_6(hash_out_valid_filter_4_6),
    .hash_out_4_7(hash_out_4_7),
    .hash_out_valid_filter_4_7(hash_out_valid_filter_4_7),
    .hash_out_5_0(hash_out_5_0),
    .hash_out_valid_filter_5_0(hash_out_valid_filter_5_0),
    .hash_out_5_1(hash_out_5_1),
    .hash_out_valid_filter_5_1(hash_out_valid_filter_5_1),
    .hash_out_5_2(hash_out_5_2),
    .hash_out_valid_filter_5_2(hash_out_valid_filter_5_2),
    .hash_out_5_3(hash_out_5_3),
    .hash_out_valid_filter_5_3(hash_out_valid_filter_5_3),
    .hash_out_5_4(hash_out_5_4),
    .hash_out_valid_filter_5_4(hash_out_valid_filter_5_4),
    .hash_out_5_5(hash_out_5_5),
    .hash_out_valid_filter_5_5(hash_out_valid_filter_5_5),
    .hash_out_5_6(hash_out_5_6),
    .hash_out_valid_filter_5_6(hash_out_valid_filter_5_6),
    .hash_out_5_7(hash_out_5_7),
    .hash_out_valid_filter_5_7(hash_out_valid_filter_5_7),
    .hash_out_6_0(hash_out_6_0),
    .hash_out_valid_filter_6_0(hash_out_valid_filter_6_0),
    .hash_out_6_1(hash_out_6_1),
    .hash_out_valid_filter_6_1(hash_out_valid_filter_6_1),
    .hash_out_6_2(hash_out_6_2),
    .hash_out_valid_filter_6_2(hash_out_valid_filter_6_2),
    .hash_out_6_3(hash_out_6_3),
    .hash_out_valid_filter_6_3(hash_out_valid_filter_6_3),
    .hash_out_6_4(hash_out_6_4),
    .hash_out_valid_filter_6_4(hash_out_valid_filter_6_4),
    .hash_out_6_5(hash_out_6_5),
    .hash_out_valid_filter_6_5(hash_out_valid_filter_6_5),
    .hash_out_6_6(hash_out_6_6),
    .hash_out_valid_filter_6_6(hash_out_valid_filter_6_6),
    .hash_out_6_7(hash_out_6_7),
    .hash_out_valid_filter_6_7(hash_out_valid_filter_6_7),
    .hash_out_7_0(hash_out_7_0),
    .hash_out_valid_filter_7_0(hash_out_valid_filter_7_0),
    .hash_out_7_1(hash_out_7_1),
    .hash_out_valid_filter_7_1(hash_out_valid_filter_7_1),
    .hash_out_7_2(hash_out_7_2),
    .hash_out_valid_filter_7_2(hash_out_valid_filter_7_2),
    .hash_out_7_3(hash_out_7_3),
    .hash_out_valid_filter_7_3(hash_out_valid_filter_7_3),
    .hash_out_7_4(hash_out_7_4),
    .hash_out_valid_filter_7_4(hash_out_valid_filter_7_4),
    .hash_out_7_5(hash_out_7_5),
    .hash_out_valid_filter_7_5(hash_out_valid_filter_7_5),
    .hash_out_7_6(hash_out_7_6),
    .hash_out_valid_filter_7_6(hash_out_valid_filter_7_6),
    .hash_out_7_7(hash_out_7_7),
    .hash_out_valid_filter_7_7(hash_out_valid_filter_7_7),
    .in_data(in_data_r2),
    .in_valid(in_valid_r2),
    .init(init_r2),
    .in_last(in_last_r2),
    .in_strb(in_strb_r2),
    .out_new_pkt(out_new_pkt)
);

//RuleID reduction logic
backend back(
    .clk(clk),
    .rst(rst),
    .din_0_0(din_0_0_r2),
    .din_valid_0_0(din_valid_0_0_r2),
    .din_almost_full_0_0(din_almost_full_0_0),
    .din_0_1(din_0_1_r2),
    .din_valid_0_1(din_valid_0_1_r2),
    .din_almost_full_0_1(din_almost_full_0_1),
    .din_0_2(din_0_2_r2),
    .din_valid_0_2(din_valid_0_2_r2),
    .din_almost_full_0_2(din_almost_full_0_2),
    .din_0_3(din_0_3_r2),
    .din_valid_0_3(din_valid_0_3_r2),
    .din_almost_full_0_3(din_almost_full_0_3),
    .din_0_4(din_0_4_r2),
    .din_valid_0_4(din_valid_0_4_r2),
    .din_almost_full_0_4(din_almost_full_0_4),
    .din_0_5(din_0_5_r2),
    .din_valid_0_5(din_valid_0_5_r2),
    .din_almost_full_0_5(din_almost_full_0_5),
    .din_0_6(din_0_6_r2),
    .din_valid_0_6(din_valid_0_6_r2),
    .din_almost_full_0_6(din_almost_full_0_6),
    .din_0_7(din_0_7_r2),
    .din_valid_0_7(din_valid_0_7_r2),
    .din_almost_full_0_7(din_almost_full_0_7),
    .din_0_8(din_0_8_r2),
    .din_valid_0_8(din_valid_0_8_r2),
    .din_almost_full_0_8(din_almost_full_0_8),
    .din_0_9(din_0_9_r2),
    .din_valid_0_9(din_valid_0_9_r2),
    .din_almost_full_0_9(din_almost_full_0_9),
    .din_0_10(din_0_10_r2),
    .din_valid_0_10(din_valid_0_10_r2),
    .din_almost_full_0_10(din_almost_full_0_10),
    .din_0_11(din_0_11_r2),
    .din_valid_0_11(din_valid_0_11_r2),
    .din_almost_full_0_11(din_almost_full_0_11),
    .din_0_12(din_0_12_r2),
    .din_valid_0_12(din_valid_0_12_r2),
    .din_almost_full_0_12(din_almost_full_0_12),
    .din_0_13(din_0_13_r2),
    .din_valid_0_13(din_valid_0_13_r2),
    .din_almost_full_0_13(din_almost_full_0_13),
    .din_0_14(din_0_14_r2),
    .din_valid_0_14(din_valid_0_14_r2),
    .din_almost_full_0_14(din_almost_full_0_14),
    .din_0_15(din_0_15_r2),
    .din_valid_0_15(din_valid_0_15_r2),
    .din_almost_full_0_15(din_almost_full_0_15),
    .din_0_16(din_0_16_r2),
    .din_valid_0_16(din_valid_0_16_r2),
    .din_almost_full_0_16(din_almost_full_0_16),
    .din_0_17(din_0_17_r2),
    .din_valid_0_17(din_valid_0_17_r2),
    .din_almost_full_0_17(din_almost_full_0_17),
    .din_0_18(din_0_18_r2),
    .din_valid_0_18(din_valid_0_18_r2),
    .din_almost_full_0_18(din_almost_full_0_18),
    .din_0_19(din_0_19_r2),
    .din_valid_0_19(din_valid_0_19_r2),
    .din_almost_full_0_19(din_almost_full_0_19),
    .din_0_20(din_0_20_r2),
    .din_valid_0_20(din_valid_0_20_r2),
    .din_almost_full_0_20(din_almost_full_0_20),
    .din_0_21(din_0_21_r2),
    .din_valid_0_21(din_valid_0_21_r2),
    .din_almost_full_0_21(din_almost_full_0_21),
    .din_0_22(din_0_22_r2),
    .din_valid_0_22(din_valid_0_22_r2),
    .din_almost_full_0_22(din_almost_full_0_22),
    .din_0_23(din_0_23_r2),
    .din_valid_0_23(din_valid_0_23_r2),
    .din_almost_full_0_23(din_almost_full_0_23),
    .din_0_24(din_0_24_r2),
    .din_valid_0_24(din_valid_0_24_r2),
    .din_almost_full_0_24(din_almost_full_0_24),
    .din_0_25(din_0_25_r2),
    .din_valid_0_25(din_valid_0_25_r2),
    .din_almost_full_0_25(din_almost_full_0_25),
    .din_0_26(din_0_26_r2),
    .din_valid_0_26(din_valid_0_26_r2),
    .din_almost_full_0_26(din_almost_full_0_26),
    .din_0_27(din_0_27_r2),
    .din_valid_0_27(din_valid_0_27_r2),
    .din_almost_full_0_27(din_almost_full_0_27),
    .din_0_28(din_0_28_r2),
    .din_valid_0_28(din_valid_0_28_r2),
    .din_almost_full_0_28(din_almost_full_0_28),
    .din_0_29(din_0_29_r2),
    .din_valid_0_29(din_valid_0_29_r2),
    .din_almost_full_0_29(din_almost_full_0_29),
    .din_0_30(din_0_30_r2),
    .din_valid_0_30(din_valid_0_30_r2),
    .din_almost_full_0_30(din_almost_full_0_30),
    .din_0_31(din_0_31_r2),
    .din_valid_0_31(din_valid_0_31_r2),
    .din_almost_full_0_31(din_almost_full_0_31),
    .din_1_0(din_1_0_r2),
    .din_valid_1_0(din_valid_1_0_r2),
    .din_almost_full_1_0(din_almost_full_1_0),
    .din_1_1(din_1_1_r2),
    .din_valid_1_1(din_valid_1_1_r2),
    .din_almost_full_1_1(din_almost_full_1_1),
    .din_1_2(din_1_2_r2),
    .din_valid_1_2(din_valid_1_2_r2),
    .din_almost_full_1_2(din_almost_full_1_2),
    .din_1_3(din_1_3_r2),
    .din_valid_1_3(din_valid_1_3_r2),
    .din_almost_full_1_3(din_almost_full_1_3),
    .din_1_4(din_1_4_r2),
    .din_valid_1_4(din_valid_1_4_r2),
    .din_almost_full_1_4(din_almost_full_1_4),
    .din_1_5(din_1_5_r2),
    .din_valid_1_5(din_valid_1_5_r2),
    .din_almost_full_1_5(din_almost_full_1_5),
    .din_1_6(din_1_6_r2),
    .din_valid_1_6(din_valid_1_6_r2),
    .din_almost_full_1_6(din_almost_full_1_6),
    .din_1_7(din_1_7_r2),
    .din_valid_1_7(din_valid_1_7_r2),
    .din_almost_full_1_7(din_almost_full_1_7),
    .din_1_8(din_1_8_r2),
    .din_valid_1_8(din_valid_1_8_r2),
    .din_almost_full_1_8(din_almost_full_1_8),
    .din_1_9(din_1_9_r2),
    .din_valid_1_9(din_valid_1_9_r2),
    .din_almost_full_1_9(din_almost_full_1_9),
    .din_1_10(din_1_10_r2),
    .din_valid_1_10(din_valid_1_10_r2),
    .din_almost_full_1_10(din_almost_full_1_10),
    .din_1_11(din_1_11_r2),
    .din_valid_1_11(din_valid_1_11_r2),
    .din_almost_full_1_11(din_almost_full_1_11),
    .din_1_12(din_1_12_r2),
    .din_valid_1_12(din_valid_1_12_r2),
    .din_almost_full_1_12(din_almost_full_1_12),
    .din_1_13(din_1_13_r2),
    .din_valid_1_13(din_valid_1_13_r2),
    .din_almost_full_1_13(din_almost_full_1_13),
    .din_1_14(din_1_14_r2),
    .din_valid_1_14(din_valid_1_14_r2),
    .din_almost_full_1_14(din_almost_full_1_14),
    .din_1_15(din_1_15_r2),
    .din_valid_1_15(din_valid_1_15_r2),
    .din_almost_full_1_15(din_almost_full_1_15),
    .din_1_16(din_1_16_r2),
    .din_valid_1_16(din_valid_1_16_r2),
    .din_almost_full_1_16(din_almost_full_1_16),
    .din_1_17(din_1_17_r2),
    .din_valid_1_17(din_valid_1_17_r2),
    .din_almost_full_1_17(din_almost_full_1_17),
    .din_1_18(din_1_18_r2),
    .din_valid_1_18(din_valid_1_18_r2),
    .din_almost_full_1_18(din_almost_full_1_18),
    .din_1_19(din_1_19_r2),
    .din_valid_1_19(din_valid_1_19_r2),
    .din_almost_full_1_19(din_almost_full_1_19),
    .din_1_20(din_1_20_r2),
    .din_valid_1_20(din_valid_1_20_r2),
    .din_almost_full_1_20(din_almost_full_1_20),
    .din_1_21(din_1_21_r2),
    .din_valid_1_21(din_valid_1_21_r2),
    .din_almost_full_1_21(din_almost_full_1_21),
    .din_1_22(din_1_22_r2),
    .din_valid_1_22(din_valid_1_22_r2),
    .din_almost_full_1_22(din_almost_full_1_22),
    .din_1_23(din_1_23_r2),
    .din_valid_1_23(din_valid_1_23_r2),
    .din_almost_full_1_23(din_almost_full_1_23),
    .din_1_24(din_1_24_r2),
    .din_valid_1_24(din_valid_1_24_r2),
    .din_almost_full_1_24(din_almost_full_1_24),
    .din_1_25(din_1_25_r2),
    .din_valid_1_25(din_valid_1_25_r2),
    .din_almost_full_1_25(din_almost_full_1_25),
    .din_1_26(din_1_26_r2),
    .din_valid_1_26(din_valid_1_26_r2),
    .din_almost_full_1_26(din_almost_full_1_26),
    .din_1_27(din_1_27_r2),
    .din_valid_1_27(din_valid_1_27_r2),
    .din_almost_full_1_27(din_almost_full_1_27),
    .din_1_28(din_1_28_r2),
    .din_valid_1_28(din_valid_1_28_r2),
    .din_almost_full_1_28(din_almost_full_1_28),
    .din_1_29(din_1_29_r2),
    .din_valid_1_29(din_valid_1_29_r2),
    .din_almost_full_1_29(din_almost_full_1_29),
    .din_1_30(din_1_30_r2),
    .din_valid_1_30(din_valid_1_30_r2),
    .din_almost_full_1_30(din_almost_full_1_30),
    .din_1_31(din_1_31_r2),
    .din_valid_1_31(din_valid_1_31_r2),
    .din_almost_full_1_31(din_almost_full_1_31),
    .din_2_0(din_2_0_r2),
    .din_valid_2_0(din_valid_2_0_r2),
    .din_almost_full_2_0(din_almost_full_2_0),
    .din_2_1(din_2_1_r2),
    .din_valid_2_1(din_valid_2_1_r2),
    .din_almost_full_2_1(din_almost_full_2_1),
    .din_2_2(din_2_2_r2),
    .din_valid_2_2(din_valid_2_2_r2),
    .din_almost_full_2_2(din_almost_full_2_2),
    .din_2_3(din_2_3_r2),
    .din_valid_2_3(din_valid_2_3_r2),
    .din_almost_full_2_3(din_almost_full_2_3),
    .din_2_4(din_2_4_r2),
    .din_valid_2_4(din_valid_2_4_r2),
    .din_almost_full_2_4(din_almost_full_2_4),
    .din_2_5(din_2_5_r2),
    .din_valid_2_5(din_valid_2_5_r2),
    .din_almost_full_2_5(din_almost_full_2_5),
    .din_2_6(din_2_6_r2),
    .din_valid_2_6(din_valid_2_6_r2),
    .din_almost_full_2_6(din_almost_full_2_6),
    .din_2_7(din_2_7_r2),
    .din_valid_2_7(din_valid_2_7_r2),
    .din_almost_full_2_7(din_almost_full_2_7),
    .din_2_8(din_2_8_r2),
    .din_valid_2_8(din_valid_2_8_r2),
    .din_almost_full_2_8(din_almost_full_2_8),
    .din_2_9(din_2_9_r2),
    .din_valid_2_9(din_valid_2_9_r2),
    .din_almost_full_2_9(din_almost_full_2_9),
    .din_2_10(din_2_10_r2),
    .din_valid_2_10(din_valid_2_10_r2),
    .din_almost_full_2_10(din_almost_full_2_10),
    .din_2_11(din_2_11_r2),
    .din_valid_2_11(din_valid_2_11_r2),
    .din_almost_full_2_11(din_almost_full_2_11),
    .din_2_12(din_2_12_r2),
    .din_valid_2_12(din_valid_2_12_r2),
    .din_almost_full_2_12(din_almost_full_2_12),
    .din_2_13(din_2_13_r2),
    .din_valid_2_13(din_valid_2_13_r2),
    .din_almost_full_2_13(din_almost_full_2_13),
    .din_2_14(din_2_14_r2),
    .din_valid_2_14(din_valid_2_14_r2),
    .din_almost_full_2_14(din_almost_full_2_14),
    .din_2_15(din_2_15_r2),
    .din_valid_2_15(din_valid_2_15_r2),
    .din_almost_full_2_15(din_almost_full_2_15),
    .din_2_16(din_2_16_r2),
    .din_valid_2_16(din_valid_2_16_r2),
    .din_almost_full_2_16(din_almost_full_2_16),
    .din_2_17(din_2_17_r2),
    .din_valid_2_17(din_valid_2_17_r2),
    .din_almost_full_2_17(din_almost_full_2_17),
    .din_2_18(din_2_18_r2),
    .din_valid_2_18(din_valid_2_18_r2),
    .din_almost_full_2_18(din_almost_full_2_18),
    .din_2_19(din_2_19_r2),
    .din_valid_2_19(din_valid_2_19_r2),
    .din_almost_full_2_19(din_almost_full_2_19),
    .din_2_20(din_2_20_r2),
    .din_valid_2_20(din_valid_2_20_r2),
    .din_almost_full_2_20(din_almost_full_2_20),
    .din_2_21(din_2_21_r2),
    .din_valid_2_21(din_valid_2_21_r2),
    .din_almost_full_2_21(din_almost_full_2_21),
    .din_2_22(din_2_22_r2),
    .din_valid_2_22(din_valid_2_22_r2),
    .din_almost_full_2_22(din_almost_full_2_22),
    .din_2_23(din_2_23_r2),
    .din_valid_2_23(din_valid_2_23_r2),
    .din_almost_full_2_23(din_almost_full_2_23),
    .din_2_24(din_2_24_r2),
    .din_valid_2_24(din_valid_2_24_r2),
    .din_almost_full_2_24(din_almost_full_2_24),
    .din_2_25(din_2_25_r2),
    .din_valid_2_25(din_valid_2_25_r2),
    .din_almost_full_2_25(din_almost_full_2_25),
    .din_2_26(din_2_26_r2),
    .din_valid_2_26(din_valid_2_26_r2),
    .din_almost_full_2_26(din_almost_full_2_26),
    .din_2_27(din_2_27_r2),
    .din_valid_2_27(din_valid_2_27_r2),
    .din_almost_full_2_27(din_almost_full_2_27),
    .din_2_28(din_2_28_r2),
    .din_valid_2_28(din_valid_2_28_r2),
    .din_almost_full_2_28(din_almost_full_2_28),
    .din_2_29(din_2_29_r2),
    .din_valid_2_29(din_valid_2_29_r2),
    .din_almost_full_2_29(din_almost_full_2_29),
    .din_2_30(din_2_30_r2),
    .din_valid_2_30(din_valid_2_30_r2),
    .din_almost_full_2_30(din_almost_full_2_30),
    .din_2_31(din_2_31_r2),
    .din_valid_2_31(din_valid_2_31_r2),
    .din_almost_full_2_31(din_almost_full_2_31),
    .din_3_0(din_3_0_r2),
    .din_valid_3_0(din_valid_3_0_r2),
    .din_almost_full_3_0(din_almost_full_3_0),
    .din_3_1(din_3_1_r2),
    .din_valid_3_1(din_valid_3_1_r2),
    .din_almost_full_3_1(din_almost_full_3_1),
    .din_3_2(din_3_2_r2),
    .din_valid_3_2(din_valid_3_2_r2),
    .din_almost_full_3_2(din_almost_full_3_2),
    .din_3_3(din_3_3_r2),
    .din_valid_3_3(din_valid_3_3_r2),
    .din_almost_full_3_3(din_almost_full_3_3),
    .din_3_4(din_3_4_r2),
    .din_valid_3_4(din_valid_3_4_r2),
    .din_almost_full_3_4(din_almost_full_3_4),
    .din_3_5(din_3_5_r2),
    .din_valid_3_5(din_valid_3_5_r2),
    .din_almost_full_3_5(din_almost_full_3_5),
    .din_3_6(din_3_6_r2),
    .din_valid_3_6(din_valid_3_6_r2),
    .din_almost_full_3_6(din_almost_full_3_6),
    .din_3_7(din_3_7_r2),
    .din_valid_3_7(din_valid_3_7_r2),
    .din_almost_full_3_7(din_almost_full_3_7),
    .din_3_8(din_3_8_r2),
    .din_valid_3_8(din_valid_3_8_r2),
    .din_almost_full_3_8(din_almost_full_3_8),
    .din_3_9(din_3_9_r2),
    .din_valid_3_9(din_valid_3_9_r2),
    .din_almost_full_3_9(din_almost_full_3_9),
    .din_3_10(din_3_10_r2),
    .din_valid_3_10(din_valid_3_10_r2),
    .din_almost_full_3_10(din_almost_full_3_10),
    .din_3_11(din_3_11_r2),
    .din_valid_3_11(din_valid_3_11_r2),
    .din_almost_full_3_11(din_almost_full_3_11),
    .din_3_12(din_3_12_r2),
    .din_valid_3_12(din_valid_3_12_r2),
    .din_almost_full_3_12(din_almost_full_3_12),
    .din_3_13(din_3_13_r2),
    .din_valid_3_13(din_valid_3_13_r2),
    .din_almost_full_3_13(din_almost_full_3_13),
    .din_3_14(din_3_14_r2),
    .din_valid_3_14(din_valid_3_14_r2),
    .din_almost_full_3_14(din_almost_full_3_14),
    .din_3_15(din_3_15_r2),
    .din_valid_3_15(din_valid_3_15_r2),
    .din_almost_full_3_15(din_almost_full_3_15),
    .din_3_16(din_3_16_r2),
    .din_valid_3_16(din_valid_3_16_r2),
    .din_almost_full_3_16(din_almost_full_3_16),
    .din_3_17(din_3_17_r2),
    .din_valid_3_17(din_valid_3_17_r2),
    .din_almost_full_3_17(din_almost_full_3_17),
    .din_3_18(din_3_18_r2),
    .din_valid_3_18(din_valid_3_18_r2),
    .din_almost_full_3_18(din_almost_full_3_18),
    .din_3_19(din_3_19_r2),
    .din_valid_3_19(din_valid_3_19_r2),
    .din_almost_full_3_19(din_almost_full_3_19),
    .din_3_20(din_3_20_r2),
    .din_valid_3_20(din_valid_3_20_r2),
    .din_almost_full_3_20(din_almost_full_3_20),
    .din_3_21(din_3_21_r2),
    .din_valid_3_21(din_valid_3_21_r2),
    .din_almost_full_3_21(din_almost_full_3_21),
    .din_3_22(din_3_22_r2),
    .din_valid_3_22(din_valid_3_22_r2),
    .din_almost_full_3_22(din_almost_full_3_22),
    .din_3_23(din_3_23_r2),
    .din_valid_3_23(din_valid_3_23_r2),
    .din_almost_full_3_23(din_almost_full_3_23),
    .din_3_24(din_3_24_r2),
    .din_valid_3_24(din_valid_3_24_r2),
    .din_almost_full_3_24(din_almost_full_3_24),
    .din_3_25(din_3_25_r2),
    .din_valid_3_25(din_valid_3_25_r2),
    .din_almost_full_3_25(din_almost_full_3_25),
    .din_3_26(din_3_26_r2),
    .din_valid_3_26(din_valid_3_26_r2),
    .din_almost_full_3_26(din_almost_full_3_26),
    .din_3_27(din_3_27_r2),
    .din_valid_3_27(din_valid_3_27_r2),
    .din_almost_full_3_27(din_almost_full_3_27),
    .din_3_28(din_3_28_r2),
    .din_valid_3_28(din_valid_3_28_r2),
    .din_almost_full_3_28(din_almost_full_3_28),
    .din_3_29(din_3_29_r2),
    .din_valid_3_29(din_valid_3_29_r2),
    .din_almost_full_3_29(din_almost_full_3_29),
    .din_3_30(din_3_30_r2),
    .din_valid_3_30(din_valid_3_30_r2),
    .din_almost_full_3_30(din_almost_full_3_30),
    .din_3_31(din_3_31_r2),
    .din_valid_3_31(din_valid_3_31_r2),
    .din_almost_full_3_31(din_almost_full_3_31),
    .din_4_0(din_4_0_r2),
    .din_valid_4_0(din_valid_4_0_r2),
    .din_almost_full_4_0(din_almost_full_4_0),
    .din_4_1(din_4_1_r2),
    .din_valid_4_1(din_valid_4_1_r2),
    .din_almost_full_4_1(din_almost_full_4_1),
    .din_4_2(din_4_2_r2),
    .din_valid_4_2(din_valid_4_2_r2),
    .din_almost_full_4_2(din_almost_full_4_2),
    .din_4_3(din_4_3_r2),
    .din_valid_4_3(din_valid_4_3_r2),
    .din_almost_full_4_3(din_almost_full_4_3),
    .din_4_4(din_4_4_r2),
    .din_valid_4_4(din_valid_4_4_r2),
    .din_almost_full_4_4(din_almost_full_4_4),
    .din_4_5(din_4_5_r2),
    .din_valid_4_5(din_valid_4_5_r2),
    .din_almost_full_4_5(din_almost_full_4_5),
    .din_4_6(din_4_6_r2),
    .din_valid_4_6(din_valid_4_6_r2),
    .din_almost_full_4_6(din_almost_full_4_6),
    .din_4_7(din_4_7_r2),
    .din_valid_4_7(din_valid_4_7_r2),
    .din_almost_full_4_7(din_almost_full_4_7),
    .din_4_8(din_4_8_r2),
    .din_valid_4_8(din_valid_4_8_r2),
    .din_almost_full_4_8(din_almost_full_4_8),
    .din_4_9(din_4_9_r2),
    .din_valid_4_9(din_valid_4_9_r2),
    .din_almost_full_4_9(din_almost_full_4_9),
    .din_4_10(din_4_10_r2),
    .din_valid_4_10(din_valid_4_10_r2),
    .din_almost_full_4_10(din_almost_full_4_10),
    .din_4_11(din_4_11_r2),
    .din_valid_4_11(din_valid_4_11_r2),
    .din_almost_full_4_11(din_almost_full_4_11),
    .din_4_12(din_4_12_r2),
    .din_valid_4_12(din_valid_4_12_r2),
    .din_almost_full_4_12(din_almost_full_4_12),
    .din_4_13(din_4_13_r2),
    .din_valid_4_13(din_valid_4_13_r2),
    .din_almost_full_4_13(din_almost_full_4_13),
    .din_4_14(din_4_14_r2),
    .din_valid_4_14(din_valid_4_14_r2),
    .din_almost_full_4_14(din_almost_full_4_14),
    .din_4_15(din_4_15_r2),
    .din_valid_4_15(din_valid_4_15_r2),
    .din_almost_full_4_15(din_almost_full_4_15),
    .din_4_16(din_4_16_r2),
    .din_valid_4_16(din_valid_4_16_r2),
    .din_almost_full_4_16(din_almost_full_4_16),
    .din_4_17(din_4_17_r2),
    .din_valid_4_17(din_valid_4_17_r2),
    .din_almost_full_4_17(din_almost_full_4_17),
    .din_4_18(din_4_18_r2),
    .din_valid_4_18(din_valid_4_18_r2),
    .din_almost_full_4_18(din_almost_full_4_18),
    .din_4_19(din_4_19_r2),
    .din_valid_4_19(din_valid_4_19_r2),
    .din_almost_full_4_19(din_almost_full_4_19),
    .din_4_20(din_4_20_r2),
    .din_valid_4_20(din_valid_4_20_r2),
    .din_almost_full_4_20(din_almost_full_4_20),
    .din_4_21(din_4_21_r2),
    .din_valid_4_21(din_valid_4_21_r2),
    .din_almost_full_4_21(din_almost_full_4_21),
    .din_4_22(din_4_22_r2),
    .din_valid_4_22(din_valid_4_22_r2),
    .din_almost_full_4_22(din_almost_full_4_22),
    .din_4_23(din_4_23_r2),
    .din_valid_4_23(din_valid_4_23_r2),
    .din_almost_full_4_23(din_almost_full_4_23),
    .din_4_24(din_4_24_r2),
    .din_valid_4_24(din_valid_4_24_r2),
    .din_almost_full_4_24(din_almost_full_4_24),
    .din_4_25(din_4_25_r2),
    .din_valid_4_25(din_valid_4_25_r2),
    .din_almost_full_4_25(din_almost_full_4_25),
    .din_4_26(din_4_26_r2),
    .din_valid_4_26(din_valid_4_26_r2),
    .din_almost_full_4_26(din_almost_full_4_26),
    .din_4_27(din_4_27_r2),
    .din_valid_4_27(din_valid_4_27_r2),
    .din_almost_full_4_27(din_almost_full_4_27),
    .din_4_28(din_4_28_r2),
    .din_valid_4_28(din_valid_4_28_r2),
    .din_almost_full_4_28(din_almost_full_4_28),
    .din_4_29(din_4_29_r2),
    .din_valid_4_29(din_valid_4_29_r2),
    .din_almost_full_4_29(din_almost_full_4_29),
    .din_4_30(din_4_30_r2),
    .din_valid_4_30(din_valid_4_30_r2),
    .din_almost_full_4_30(din_almost_full_4_30),
    .din_4_31(din_4_31_r2),
    .din_valid_4_31(din_valid_4_31_r2),
    .din_almost_full_4_31(din_almost_full_4_31),
    .din_5_0(din_5_0_r2),
    .din_valid_5_0(din_valid_5_0_r2),
    .din_almost_full_5_0(din_almost_full_5_0),
    .din_5_1(din_5_1_r2),
    .din_valid_5_1(din_valid_5_1_r2),
    .din_almost_full_5_1(din_almost_full_5_1),
    .din_5_2(din_5_2_r2),
    .din_valid_5_2(din_valid_5_2_r2),
    .din_almost_full_5_2(din_almost_full_5_2),
    .din_5_3(din_5_3_r2),
    .din_valid_5_3(din_valid_5_3_r2),
    .din_almost_full_5_3(din_almost_full_5_3),
    .din_5_4(din_5_4_r2),
    .din_valid_5_4(din_valid_5_4_r2),
    .din_almost_full_5_4(din_almost_full_5_4),
    .din_5_5(din_5_5_r2),
    .din_valid_5_5(din_valid_5_5_r2),
    .din_almost_full_5_5(din_almost_full_5_5),
    .din_5_6(din_5_6_r2),
    .din_valid_5_6(din_valid_5_6_r2),
    .din_almost_full_5_6(din_almost_full_5_6),
    .din_5_7(din_5_7_r2),
    .din_valid_5_7(din_valid_5_7_r2),
    .din_almost_full_5_7(din_almost_full_5_7),
    .din_5_8(din_5_8_r2),
    .din_valid_5_8(din_valid_5_8_r2),
    .din_almost_full_5_8(din_almost_full_5_8),
    .din_5_9(din_5_9_r2),
    .din_valid_5_9(din_valid_5_9_r2),
    .din_almost_full_5_9(din_almost_full_5_9),
    .din_5_10(din_5_10_r2),
    .din_valid_5_10(din_valid_5_10_r2),
    .din_almost_full_5_10(din_almost_full_5_10),
    .din_5_11(din_5_11_r2),
    .din_valid_5_11(din_valid_5_11_r2),
    .din_almost_full_5_11(din_almost_full_5_11),
    .din_5_12(din_5_12_r2),
    .din_valid_5_12(din_valid_5_12_r2),
    .din_almost_full_5_12(din_almost_full_5_12),
    .din_5_13(din_5_13_r2),
    .din_valid_5_13(din_valid_5_13_r2),
    .din_almost_full_5_13(din_almost_full_5_13),
    .din_5_14(din_5_14_r2),
    .din_valid_5_14(din_valid_5_14_r2),
    .din_almost_full_5_14(din_almost_full_5_14),
    .din_5_15(din_5_15_r2),
    .din_valid_5_15(din_valid_5_15_r2),
    .din_almost_full_5_15(din_almost_full_5_15),
    .din_5_16(din_5_16_r2),
    .din_valid_5_16(din_valid_5_16_r2),
    .din_almost_full_5_16(din_almost_full_5_16),
    .din_5_17(din_5_17_r2),
    .din_valid_5_17(din_valid_5_17_r2),
    .din_almost_full_5_17(din_almost_full_5_17),
    .din_5_18(din_5_18_r2),
    .din_valid_5_18(din_valid_5_18_r2),
    .din_almost_full_5_18(din_almost_full_5_18),
    .din_5_19(din_5_19_r2),
    .din_valid_5_19(din_valid_5_19_r2),
    .din_almost_full_5_19(din_almost_full_5_19),
    .din_5_20(din_5_20_r2),
    .din_valid_5_20(din_valid_5_20_r2),
    .din_almost_full_5_20(din_almost_full_5_20),
    .din_5_21(din_5_21_r2),
    .din_valid_5_21(din_valid_5_21_r2),
    .din_almost_full_5_21(din_almost_full_5_21),
    .din_5_22(din_5_22_r2),
    .din_valid_5_22(din_valid_5_22_r2),
    .din_almost_full_5_22(din_almost_full_5_22),
    .din_5_23(din_5_23_r2),
    .din_valid_5_23(din_valid_5_23_r2),
    .din_almost_full_5_23(din_almost_full_5_23),
    .din_5_24(din_5_24_r2),
    .din_valid_5_24(din_valid_5_24_r2),
    .din_almost_full_5_24(din_almost_full_5_24),
    .din_5_25(din_5_25_r2),
    .din_valid_5_25(din_valid_5_25_r2),
    .din_almost_full_5_25(din_almost_full_5_25),
    .din_5_26(din_5_26_r2),
    .din_valid_5_26(din_valid_5_26_r2),
    .din_almost_full_5_26(din_almost_full_5_26),
    .din_5_27(din_5_27_r2),
    .din_valid_5_27(din_valid_5_27_r2),
    .din_almost_full_5_27(din_almost_full_5_27),
    .din_5_28(din_5_28_r2),
    .din_valid_5_28(din_valid_5_28_r2),
    .din_almost_full_5_28(din_almost_full_5_28),
    .din_5_29(din_5_29_r2),
    .din_valid_5_29(din_valid_5_29_r2),
    .din_almost_full_5_29(din_almost_full_5_29),
    .din_5_30(din_5_30_r2),
    .din_valid_5_30(din_valid_5_30_r2),
    .din_almost_full_5_30(din_almost_full_5_30),
    .din_5_31(din_5_31_r2),
    .din_valid_5_31(din_valid_5_31_r2),
    .din_almost_full_5_31(din_almost_full_5_31),
    .din_6_0(din_6_0_r2),
    .din_valid_6_0(din_valid_6_0_r2),
    .din_almost_full_6_0(din_almost_full_6_0),
    .din_6_1(din_6_1_r2),
    .din_valid_6_1(din_valid_6_1_r2),
    .din_almost_full_6_1(din_almost_full_6_1),
    .din_6_2(din_6_2_r2),
    .din_valid_6_2(din_valid_6_2_r2),
    .din_almost_full_6_2(din_almost_full_6_2),
    .din_6_3(din_6_3_r2),
    .din_valid_6_3(din_valid_6_3_r2),
    .din_almost_full_6_3(din_almost_full_6_3),
    .din_6_4(din_6_4_r2),
    .din_valid_6_4(din_valid_6_4_r2),
    .din_almost_full_6_4(din_almost_full_6_4),
    .din_6_5(din_6_5_r2),
    .din_valid_6_5(din_valid_6_5_r2),
    .din_almost_full_6_5(din_almost_full_6_5),
    .din_6_6(din_6_6_r2),
    .din_valid_6_6(din_valid_6_6_r2),
    .din_almost_full_6_6(din_almost_full_6_6),
    .din_6_7(din_6_7_r2),
    .din_valid_6_7(din_valid_6_7_r2),
    .din_almost_full_6_7(din_almost_full_6_7),
    .din_6_8(din_6_8_r2),
    .din_valid_6_8(din_valid_6_8_r2),
    .din_almost_full_6_8(din_almost_full_6_8),
    .din_6_9(din_6_9_r2),
    .din_valid_6_9(din_valid_6_9_r2),
    .din_almost_full_6_9(din_almost_full_6_9),
    .din_6_10(din_6_10_r2),
    .din_valid_6_10(din_valid_6_10_r2),
    .din_almost_full_6_10(din_almost_full_6_10),
    .din_6_11(din_6_11_r2),
    .din_valid_6_11(din_valid_6_11_r2),
    .din_almost_full_6_11(din_almost_full_6_11),
    .din_6_12(din_6_12_r2),
    .din_valid_6_12(din_valid_6_12_r2),
    .din_almost_full_6_12(din_almost_full_6_12),
    .din_6_13(din_6_13_r2),
    .din_valid_6_13(din_valid_6_13_r2),
    .din_almost_full_6_13(din_almost_full_6_13),
    .din_6_14(din_6_14_r2),
    .din_valid_6_14(din_valid_6_14_r2),
    .din_almost_full_6_14(din_almost_full_6_14),
    .din_6_15(din_6_15_r2),
    .din_valid_6_15(din_valid_6_15_r2),
    .din_almost_full_6_15(din_almost_full_6_15),
    .din_6_16(din_6_16_r2),
    .din_valid_6_16(din_valid_6_16_r2),
    .din_almost_full_6_16(din_almost_full_6_16),
    .din_6_17(din_6_17_r2),
    .din_valid_6_17(din_valid_6_17_r2),
    .din_almost_full_6_17(din_almost_full_6_17),
    .din_6_18(din_6_18_r2),
    .din_valid_6_18(din_valid_6_18_r2),
    .din_almost_full_6_18(din_almost_full_6_18),
    .din_6_19(din_6_19_r2),
    .din_valid_6_19(din_valid_6_19_r2),
    .din_almost_full_6_19(din_almost_full_6_19),
    .din_6_20(din_6_20_r2),
    .din_valid_6_20(din_valid_6_20_r2),
    .din_almost_full_6_20(din_almost_full_6_20),
    .din_6_21(din_6_21_r2),
    .din_valid_6_21(din_valid_6_21_r2),
    .din_almost_full_6_21(din_almost_full_6_21),
    .din_6_22(din_6_22_r2),
    .din_valid_6_22(din_valid_6_22_r2),
    .din_almost_full_6_22(din_almost_full_6_22),
    .din_6_23(din_6_23_r2),
    .din_valid_6_23(din_valid_6_23_r2),
    .din_almost_full_6_23(din_almost_full_6_23),
    .din_6_24(din_6_24_r2),
    .din_valid_6_24(din_valid_6_24_r2),
    .din_almost_full_6_24(din_almost_full_6_24),
    .din_6_25(din_6_25_r2),
    .din_valid_6_25(din_valid_6_25_r2),
    .din_almost_full_6_25(din_almost_full_6_25),
    .din_6_26(din_6_26_r2),
    .din_valid_6_26(din_valid_6_26_r2),
    .din_almost_full_6_26(din_almost_full_6_26),
    .din_6_27(din_6_27_r2),
    .din_valid_6_27(din_valid_6_27_r2),
    .din_almost_full_6_27(din_almost_full_6_27),
    .din_6_28(din_6_28_r2),
    .din_valid_6_28(din_valid_6_28_r2),
    .din_almost_full_6_28(din_almost_full_6_28),
    .din_6_29(din_6_29_r2),
    .din_valid_6_29(din_valid_6_29_r2),
    .din_almost_full_6_29(din_almost_full_6_29),
    .din_6_30(din_6_30_r2),
    .din_valid_6_30(din_valid_6_30_r2),
    .din_almost_full_6_30(din_almost_full_6_30),
    .din_6_31(din_6_31_r2),
    .din_valid_6_31(din_valid_6_31_r2),
    .din_almost_full_6_31(din_almost_full_6_31),
    .din_7_0(din_7_0_r2),
    .din_valid_7_0(din_valid_7_0_r2),
    .din_almost_full_7_0(din_almost_full_7_0),
    .din_7_1(din_7_1_r2),
    .din_valid_7_1(din_valid_7_1_r2),
    .din_almost_full_7_1(din_almost_full_7_1),
    .din_7_2(din_7_2_r2),
    .din_valid_7_2(din_valid_7_2_r2),
    .din_almost_full_7_2(din_almost_full_7_2),
    .din_7_3(din_7_3_r2),
    .din_valid_7_3(din_valid_7_3_r2),
    .din_almost_full_7_3(din_almost_full_7_3),
    .din_7_4(din_7_4_r2),
    .din_valid_7_4(din_valid_7_4_r2),
    .din_almost_full_7_4(din_almost_full_7_4),
    .din_7_5(din_7_5_r2),
    .din_valid_7_5(din_valid_7_5_r2),
    .din_almost_full_7_5(din_almost_full_7_5),
    .din_7_6(din_7_6_r2),
    .din_valid_7_6(din_valid_7_6_r2),
    .din_almost_full_7_6(din_almost_full_7_6),
    .din_7_7(din_7_7_r2),
    .din_valid_7_7(din_valid_7_7_r2),
    .din_almost_full_7_7(din_almost_full_7_7),
    .din_7_8(din_7_8_r2),
    .din_valid_7_8(din_valid_7_8_r2),
    .din_almost_full_7_8(din_almost_full_7_8),
    .din_7_9(din_7_9_r2),
    .din_valid_7_9(din_valid_7_9_r2),
    .din_almost_full_7_9(din_almost_full_7_9),
    .din_7_10(din_7_10_r2),
    .din_valid_7_10(din_valid_7_10_r2),
    .din_almost_full_7_10(din_almost_full_7_10),
    .din_7_11(din_7_11_r2),
    .din_valid_7_11(din_valid_7_11_r2),
    .din_almost_full_7_11(din_almost_full_7_11),
    .din_7_12(din_7_12_r2),
    .din_valid_7_12(din_valid_7_12_r2),
    .din_almost_full_7_12(din_almost_full_7_12),
    .din_7_13(din_7_13_r2),
    .din_valid_7_13(din_valid_7_13_r2),
    .din_almost_full_7_13(din_almost_full_7_13),
    .din_7_14(din_7_14_r2),
    .din_valid_7_14(din_valid_7_14_r2),
    .din_almost_full_7_14(din_almost_full_7_14),
    .din_7_15(din_7_15_r2),
    .din_valid_7_15(din_valid_7_15_r2),
    .din_almost_full_7_15(din_almost_full_7_15),
    .din_7_16(din_7_16_r2),
    .din_valid_7_16(din_valid_7_16_r2),
    .din_almost_full_7_16(din_almost_full_7_16),
    .din_7_17(din_7_17_r2),
    .din_valid_7_17(din_valid_7_17_r2),
    .din_almost_full_7_17(din_almost_full_7_17),
    .din_7_18(din_7_18_r2),
    .din_valid_7_18(din_valid_7_18_r2),
    .din_almost_full_7_18(din_almost_full_7_18),
    .din_7_19(din_7_19_r2),
    .din_valid_7_19(din_valid_7_19_r2),
    .din_almost_full_7_19(din_almost_full_7_19),
    .din_7_20(din_7_20_r2),
    .din_valid_7_20(din_valid_7_20_r2),
    .din_almost_full_7_20(din_almost_full_7_20),
    .din_7_21(din_7_21_r2),
    .din_valid_7_21(din_valid_7_21_r2),
    .din_almost_full_7_21(din_almost_full_7_21),
    .din_7_22(din_7_22_r2),
    .din_valid_7_22(din_valid_7_22_r2),
    .din_almost_full_7_22(din_almost_full_7_22),
    .din_7_23(din_7_23_r2),
    .din_valid_7_23(din_valid_7_23_r2),
    .din_almost_full_7_23(din_almost_full_7_23),
    .din_7_24(din_7_24_r2),
    .din_valid_7_24(din_valid_7_24_r2),
    .din_almost_full_7_24(din_almost_full_7_24),
    .din_7_25(din_7_25_r2),
    .din_valid_7_25(din_valid_7_25_r2),
    .din_almost_full_7_25(din_almost_full_7_25),
    .din_7_26(din_7_26_r2),
    .din_valid_7_26(din_valid_7_26_r2),
    .din_almost_full_7_26(din_almost_full_7_26),
    .din_7_27(din_7_27_r2),
    .din_valid_7_27(din_valid_7_27_r2),
    .din_almost_full_7_27(din_almost_full_7_27),
    .din_7_28(din_7_28_r2),
    .din_valid_7_28(din_valid_7_28_r2),
    .din_almost_full_7_28(din_almost_full_7_28),
    .din_7_29(din_7_29_r2),
    .din_valid_7_29(din_valid_7_29_r2),
    .din_almost_full_7_29(din_almost_full_7_29),
    .din_7_30(din_7_30_r2),
    .din_valid_7_30(din_valid_7_30_r2),
    .din_almost_full_7_30(din_almost_full_7_30),
    .din_7_31(din_7_31_r2),
    .din_valid_7_31(din_valid_7_31_r2),
    .din_almost_full_7_31(din_almost_full_7_31),
    .ruleID(out_data),
    .ruleID_valid(out_valid),
    .ruleID_last(out_last),
    .ruleID_almost_full(out_almost_full)
);

endmodule //top
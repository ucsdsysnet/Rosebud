`include "struct_s.sv"
module hashtable_top(clk,
	dout_0_0,dout_valid_0_0,
	dout_0_1,dout_valid_0_1,
	dout_0_2,dout_valid_0_2,
	dout_0_3,dout_valid_0_3,
	dout_0_4,dout_valid_0_4,
	dout_0_5,dout_valid_0_5,
	dout_0_6,dout_valid_0_6,
	dout_0_7,dout_valid_0_7,
	dout_0_8,dout_valid_0_8,
	dout_0_9,dout_valid_0_9,
	dout_0_10,dout_valid_0_10,
	dout_0_11,dout_valid_0_11,
	dout_0_12,dout_valid_0_12,
	dout_0_13,dout_valid_0_13,
	dout_0_14,dout_valid_0_14,
	dout_0_15,dout_valid_0_15,
	dout_0_16,dout_valid_0_16,
	dout_0_17,dout_valid_0_17,
	dout_0_18,dout_valid_0_18,
	dout_0_19,dout_valid_0_19,
	dout_0_20,dout_valid_0_20,
	dout_0_21,dout_valid_0_21,
	dout_0_22,dout_valid_0_22,
	dout_0_23,dout_valid_0_23,
	dout_0_24,dout_valid_0_24,
	dout_0_25,dout_valid_0_25,
	dout_0_26,dout_valid_0_26,
	dout_0_27,dout_valid_0_27,
	dout_0_28,dout_valid_0_28,
	dout_0_29,dout_valid_0_29,
	dout_0_30,dout_valid_0_30,
	dout_0_31,dout_valid_0_31,
	dout_1_0,dout_valid_1_0,
	dout_1_1,dout_valid_1_1,
	dout_1_2,dout_valid_1_2,
	dout_1_3,dout_valid_1_3,
	dout_1_4,dout_valid_1_4,
	dout_1_5,dout_valid_1_5,
	dout_1_6,dout_valid_1_6,
	dout_1_7,dout_valid_1_7,
	dout_1_8,dout_valid_1_8,
	dout_1_9,dout_valid_1_9,
	dout_1_10,dout_valid_1_10,
	dout_1_11,dout_valid_1_11,
	dout_1_12,dout_valid_1_12,
	dout_1_13,dout_valid_1_13,
	dout_1_14,dout_valid_1_14,
	dout_1_15,dout_valid_1_15,
	dout_1_16,dout_valid_1_16,
	dout_1_17,dout_valid_1_17,
	dout_1_18,dout_valid_1_18,
	dout_1_19,dout_valid_1_19,
	dout_1_20,dout_valid_1_20,
	dout_1_21,dout_valid_1_21,
	dout_1_22,dout_valid_1_22,
	dout_1_23,dout_valid_1_23,
	dout_1_24,dout_valid_1_24,
	dout_1_25,dout_valid_1_25,
	dout_1_26,dout_valid_1_26,
	dout_1_27,dout_valid_1_27,
	dout_1_28,dout_valid_1_28,
	dout_1_29,dout_valid_1_29,
	dout_1_30,dout_valid_1_30,
	dout_1_31,dout_valid_1_31,
	dout_2_0,dout_valid_2_0,
	dout_2_1,dout_valid_2_1,
	dout_2_2,dout_valid_2_2,
	dout_2_3,dout_valid_2_3,
	dout_2_4,dout_valid_2_4,
	dout_2_5,dout_valid_2_5,
	dout_2_6,dout_valid_2_6,
	dout_2_7,dout_valid_2_7,
	dout_2_8,dout_valid_2_8,
	dout_2_9,dout_valid_2_9,
	dout_2_10,dout_valid_2_10,
	dout_2_11,dout_valid_2_11,
	dout_2_12,dout_valid_2_12,
	dout_2_13,dout_valid_2_13,
	dout_2_14,dout_valid_2_14,
	dout_2_15,dout_valid_2_15,
	dout_2_16,dout_valid_2_16,
	dout_2_17,dout_valid_2_17,
	dout_2_18,dout_valid_2_18,
	dout_2_19,dout_valid_2_19,
	dout_2_20,dout_valid_2_20,
	dout_2_21,dout_valid_2_21,
	dout_2_22,dout_valid_2_22,
	dout_2_23,dout_valid_2_23,
	dout_2_24,dout_valid_2_24,
	dout_2_25,dout_valid_2_25,
	dout_2_26,dout_valid_2_26,
	dout_2_27,dout_valid_2_27,
	dout_2_28,dout_valid_2_28,
	dout_2_29,dout_valid_2_29,
	dout_2_30,dout_valid_2_30,
	dout_2_31,dout_valid_2_31,
	dout_3_0,dout_valid_3_0,
	dout_3_1,dout_valid_3_1,
	dout_3_2,dout_valid_3_2,
	dout_3_3,dout_valid_3_3,
	dout_3_4,dout_valid_3_4,
	dout_3_5,dout_valid_3_5,
	dout_3_6,dout_valid_3_6,
	dout_3_7,dout_valid_3_7,
	dout_3_8,dout_valid_3_8,
	dout_3_9,dout_valid_3_9,
	dout_3_10,dout_valid_3_10,
	dout_3_11,dout_valid_3_11,
	dout_3_12,dout_valid_3_12,
	dout_3_13,dout_valid_3_13,
	dout_3_14,dout_valid_3_14,
	dout_3_15,dout_valid_3_15,
	dout_3_16,dout_valid_3_16,
	dout_3_17,dout_valid_3_17,
	dout_3_18,dout_valid_3_18,
	dout_3_19,dout_valid_3_19,
	dout_3_20,dout_valid_3_20,
	dout_3_21,dout_valid_3_21,
	dout_3_22,dout_valid_3_22,
	dout_3_23,dout_valid_3_23,
	dout_3_24,dout_valid_3_24,
	dout_3_25,dout_valid_3_25,
	dout_3_26,dout_valid_3_26,
	dout_3_27,dout_valid_3_27,
	dout_3_28,dout_valid_3_28,
	dout_3_29,dout_valid_3_29,
	dout_3_30,dout_valid_3_30,
	dout_3_31,dout_valid_3_31,
	dout_4_0,dout_valid_4_0,
	dout_4_1,dout_valid_4_1,
	dout_4_2,dout_valid_4_2,
	dout_4_3,dout_valid_4_3,
	dout_4_4,dout_valid_4_4,
	dout_4_5,dout_valid_4_5,
	dout_4_6,dout_valid_4_6,
	dout_4_7,dout_valid_4_7,
	dout_4_8,dout_valid_4_8,
	dout_4_9,dout_valid_4_9,
	dout_4_10,dout_valid_4_10,
	dout_4_11,dout_valid_4_11,
	dout_4_12,dout_valid_4_12,
	dout_4_13,dout_valid_4_13,
	dout_4_14,dout_valid_4_14,
	dout_4_15,dout_valid_4_15,
	dout_4_16,dout_valid_4_16,
	dout_4_17,dout_valid_4_17,
	dout_4_18,dout_valid_4_18,
	dout_4_19,dout_valid_4_19,
	dout_4_20,dout_valid_4_20,
	dout_4_21,dout_valid_4_21,
	dout_4_22,dout_valid_4_22,
	dout_4_23,dout_valid_4_23,
	dout_4_24,dout_valid_4_24,
	dout_4_25,dout_valid_4_25,
	dout_4_26,dout_valid_4_26,
	dout_4_27,dout_valid_4_27,
	dout_4_28,dout_valid_4_28,
	dout_4_29,dout_valid_4_29,
	dout_4_30,dout_valid_4_30,
	dout_4_31,dout_valid_4_31,
	dout_5_0,dout_valid_5_0,
	dout_5_1,dout_valid_5_1,
	dout_5_2,dout_valid_5_2,
	dout_5_3,dout_valid_5_3,
	dout_5_4,dout_valid_5_4,
	dout_5_5,dout_valid_5_5,
	dout_5_6,dout_valid_5_6,
	dout_5_7,dout_valid_5_7,
	dout_5_8,dout_valid_5_8,
	dout_5_9,dout_valid_5_9,
	dout_5_10,dout_valid_5_10,
	dout_5_11,dout_valid_5_11,
	dout_5_12,dout_valid_5_12,
	dout_5_13,dout_valid_5_13,
	dout_5_14,dout_valid_5_14,
	dout_5_15,dout_valid_5_15,
	dout_5_16,dout_valid_5_16,
	dout_5_17,dout_valid_5_17,
	dout_5_18,dout_valid_5_18,
	dout_5_19,dout_valid_5_19,
	dout_5_20,dout_valid_5_20,
	dout_5_21,dout_valid_5_21,
	dout_5_22,dout_valid_5_22,
	dout_5_23,dout_valid_5_23,
	dout_5_24,dout_valid_5_24,
	dout_5_25,dout_valid_5_25,
	dout_5_26,dout_valid_5_26,
	dout_5_27,dout_valid_5_27,
	dout_5_28,dout_valid_5_28,
	dout_5_29,dout_valid_5_29,
	dout_5_30,dout_valid_5_30,
	dout_5_31,dout_valid_5_31,
	dout_6_0,dout_valid_6_0,
	dout_6_1,dout_valid_6_1,
	dout_6_2,dout_valid_6_2,
	dout_6_3,dout_valid_6_3,
	dout_6_4,dout_valid_6_4,
	dout_6_5,dout_valid_6_5,
	dout_6_6,dout_valid_6_6,
	dout_6_7,dout_valid_6_7,
	dout_6_8,dout_valid_6_8,
	dout_6_9,dout_valid_6_9,
	dout_6_10,dout_valid_6_10,
	dout_6_11,dout_valid_6_11,
	dout_6_12,dout_valid_6_12,
	dout_6_13,dout_valid_6_13,
	dout_6_14,dout_valid_6_14,
	dout_6_15,dout_valid_6_15,
	dout_6_16,dout_valid_6_16,
	dout_6_17,dout_valid_6_17,
	dout_6_18,dout_valid_6_18,
	dout_6_19,dout_valid_6_19,
	dout_6_20,dout_valid_6_20,
	dout_6_21,dout_valid_6_21,
	dout_6_22,dout_valid_6_22,
	dout_6_23,dout_valid_6_23,
	dout_6_24,dout_valid_6_24,
	dout_6_25,dout_valid_6_25,
	dout_6_26,dout_valid_6_26,
	dout_6_27,dout_valid_6_27,
	dout_6_28,dout_valid_6_28,
	dout_6_29,dout_valid_6_29,
	dout_6_30,dout_valid_6_30,
	dout_6_31,dout_valid_6_31,
	dout_7_0,dout_valid_7_0,
	dout_7_1,dout_valid_7_1,
	dout_7_2,dout_valid_7_2,
	dout_7_3,dout_valid_7_3,
	dout_7_4,dout_valid_7_4,
	dout_7_5,dout_valid_7_5,
	dout_7_6,dout_valid_7_6,
	dout_7_7,dout_valid_7_7,
	dout_7_8,dout_valid_7_8,
	dout_7_9,dout_valid_7_9,
	dout_7_10,dout_valid_7_10,
	dout_7_11,dout_valid_7_11,
	dout_7_12,dout_valid_7_12,
	dout_7_13,dout_valid_7_13,
	dout_7_14,dout_valid_7_14,
	dout_7_15,dout_valid_7_15,
	dout_7_16,dout_valid_7_16,
	dout_7_17,dout_valid_7_17,
	dout_7_18,dout_valid_7_18,
	dout_7_19,dout_valid_7_19,
	dout_7_20,dout_valid_7_20,
	dout_7_21,dout_valid_7_21,
	dout_7_22,dout_valid_7_22,
	dout_7_23,dout_valid_7_23,
	dout_7_24,dout_valid_7_24,
	dout_7_25,dout_valid_7_25,
	dout_7_26,dout_valid_7_26,
	dout_7_27,dout_valid_7_27,
	dout_7_28,dout_valid_7_28,
	dout_7_29,dout_valid_7_29,
	dout_7_30,dout_valid_7_30,
	dout_7_31,dout_valid_7_31,
    din,din_valid
);

input clk;
input [255:0] din;
input din_valid;
output wire [RID_WIDTH-1:0] dout_0_0;
output wire dout_valid_0_0;
output wire [RID_WIDTH-1:0] dout_0_1;
output wire dout_valid_0_1;
output wire [RID_WIDTH-1:0] dout_0_2;
output wire dout_valid_0_2;
output wire [RID_WIDTH-1:0] dout_0_3;
output wire dout_valid_0_3;
output wire [RID_WIDTH-1:0] dout_0_4;
output wire dout_valid_0_4;
output wire [RID_WIDTH-1:0] dout_0_5;
output wire dout_valid_0_5;
output wire [RID_WIDTH-1:0] dout_0_6;
output wire dout_valid_0_6;
output wire [RID_WIDTH-1:0] dout_0_7;
output wire dout_valid_0_7;
output wire [RID_WIDTH-1:0] dout_0_8;
output wire dout_valid_0_8;
output wire [RID_WIDTH-1:0] dout_0_9;
output wire dout_valid_0_9;
output wire [RID_WIDTH-1:0] dout_0_10;
output wire dout_valid_0_10;
output wire [RID_WIDTH-1:0] dout_0_11;
output wire dout_valid_0_11;
output wire [RID_WIDTH-1:0] dout_0_12;
output wire dout_valid_0_12;
output wire [RID_WIDTH-1:0] dout_0_13;
output wire dout_valid_0_13;
output wire [RID_WIDTH-1:0] dout_0_14;
output wire dout_valid_0_14;
output wire [RID_WIDTH-1:0] dout_0_15;
output wire dout_valid_0_15;
output wire [RID_WIDTH-1:0] dout_0_16;
output wire dout_valid_0_16;
output wire [RID_WIDTH-1:0] dout_0_17;
output wire dout_valid_0_17;
output wire [RID_WIDTH-1:0] dout_0_18;
output wire dout_valid_0_18;
output wire [RID_WIDTH-1:0] dout_0_19;
output wire dout_valid_0_19;
output wire [RID_WIDTH-1:0] dout_0_20;
output wire dout_valid_0_20;
output wire [RID_WIDTH-1:0] dout_0_21;
output wire dout_valid_0_21;
output wire [RID_WIDTH-1:0] dout_0_22;
output wire dout_valid_0_22;
output wire [RID_WIDTH-1:0] dout_0_23;
output wire dout_valid_0_23;
output wire [RID_WIDTH-1:0] dout_0_24;
output wire dout_valid_0_24;
output wire [RID_WIDTH-1:0] dout_0_25;
output wire dout_valid_0_25;
output wire [RID_WIDTH-1:0] dout_0_26;
output wire dout_valid_0_26;
output wire [RID_WIDTH-1:0] dout_0_27;
output wire dout_valid_0_27;
output wire [RID_WIDTH-1:0] dout_0_28;
output wire dout_valid_0_28;
output wire [RID_WIDTH-1:0] dout_0_29;
output wire dout_valid_0_29;
output wire [RID_WIDTH-1:0] dout_0_30;
output wire dout_valid_0_30;
output wire [RID_WIDTH-1:0] dout_0_31;
output wire dout_valid_0_31;
output wire [RID_WIDTH-1:0] dout_1_0;
output wire dout_valid_1_0;
output wire [RID_WIDTH-1:0] dout_1_1;
output wire dout_valid_1_1;
output wire [RID_WIDTH-1:0] dout_1_2;
output wire dout_valid_1_2;
output wire [RID_WIDTH-1:0] dout_1_3;
output wire dout_valid_1_3;
output wire [RID_WIDTH-1:0] dout_1_4;
output wire dout_valid_1_4;
output wire [RID_WIDTH-1:0] dout_1_5;
output wire dout_valid_1_5;
output wire [RID_WIDTH-1:0] dout_1_6;
output wire dout_valid_1_6;
output wire [RID_WIDTH-1:0] dout_1_7;
output wire dout_valid_1_7;
output wire [RID_WIDTH-1:0] dout_1_8;
output wire dout_valid_1_8;
output wire [RID_WIDTH-1:0] dout_1_9;
output wire dout_valid_1_9;
output wire [RID_WIDTH-1:0] dout_1_10;
output wire dout_valid_1_10;
output wire [RID_WIDTH-1:0] dout_1_11;
output wire dout_valid_1_11;
output wire [RID_WIDTH-1:0] dout_1_12;
output wire dout_valid_1_12;
output wire [RID_WIDTH-1:0] dout_1_13;
output wire dout_valid_1_13;
output wire [RID_WIDTH-1:0] dout_1_14;
output wire dout_valid_1_14;
output wire [RID_WIDTH-1:0] dout_1_15;
output wire dout_valid_1_15;
output wire [RID_WIDTH-1:0] dout_1_16;
output wire dout_valid_1_16;
output wire [RID_WIDTH-1:0] dout_1_17;
output wire dout_valid_1_17;
output wire [RID_WIDTH-1:0] dout_1_18;
output wire dout_valid_1_18;
output wire [RID_WIDTH-1:0] dout_1_19;
output wire dout_valid_1_19;
output wire [RID_WIDTH-1:0] dout_1_20;
output wire dout_valid_1_20;
output wire [RID_WIDTH-1:0] dout_1_21;
output wire dout_valid_1_21;
output wire [RID_WIDTH-1:0] dout_1_22;
output wire dout_valid_1_22;
output wire [RID_WIDTH-1:0] dout_1_23;
output wire dout_valid_1_23;
output wire [RID_WIDTH-1:0] dout_1_24;
output wire dout_valid_1_24;
output wire [RID_WIDTH-1:0] dout_1_25;
output wire dout_valid_1_25;
output wire [RID_WIDTH-1:0] dout_1_26;
output wire dout_valid_1_26;
output wire [RID_WIDTH-1:0] dout_1_27;
output wire dout_valid_1_27;
output wire [RID_WIDTH-1:0] dout_1_28;
output wire dout_valid_1_28;
output wire [RID_WIDTH-1:0] dout_1_29;
output wire dout_valid_1_29;
output wire [RID_WIDTH-1:0] dout_1_30;
output wire dout_valid_1_30;
output wire [RID_WIDTH-1:0] dout_1_31;
output wire dout_valid_1_31;
output wire [RID_WIDTH-1:0] dout_2_0;
output wire dout_valid_2_0;
output wire [RID_WIDTH-1:0] dout_2_1;
output wire dout_valid_2_1;
output wire [RID_WIDTH-1:0] dout_2_2;
output wire dout_valid_2_2;
output wire [RID_WIDTH-1:0] dout_2_3;
output wire dout_valid_2_3;
output wire [RID_WIDTH-1:0] dout_2_4;
output wire dout_valid_2_4;
output wire [RID_WIDTH-1:0] dout_2_5;
output wire dout_valid_2_5;
output wire [RID_WIDTH-1:0] dout_2_6;
output wire dout_valid_2_6;
output wire [RID_WIDTH-1:0] dout_2_7;
output wire dout_valid_2_7;
output wire [RID_WIDTH-1:0] dout_2_8;
output wire dout_valid_2_8;
output wire [RID_WIDTH-1:0] dout_2_9;
output wire dout_valid_2_9;
output wire [RID_WIDTH-1:0] dout_2_10;
output wire dout_valid_2_10;
output wire [RID_WIDTH-1:0] dout_2_11;
output wire dout_valid_2_11;
output wire [RID_WIDTH-1:0] dout_2_12;
output wire dout_valid_2_12;
output wire [RID_WIDTH-1:0] dout_2_13;
output wire dout_valid_2_13;
output wire [RID_WIDTH-1:0] dout_2_14;
output wire dout_valid_2_14;
output wire [RID_WIDTH-1:0] dout_2_15;
output wire dout_valid_2_15;
output wire [RID_WIDTH-1:0] dout_2_16;
output wire dout_valid_2_16;
output wire [RID_WIDTH-1:0] dout_2_17;
output wire dout_valid_2_17;
output wire [RID_WIDTH-1:0] dout_2_18;
output wire dout_valid_2_18;
output wire [RID_WIDTH-1:0] dout_2_19;
output wire dout_valid_2_19;
output wire [RID_WIDTH-1:0] dout_2_20;
output wire dout_valid_2_20;
output wire [RID_WIDTH-1:0] dout_2_21;
output wire dout_valid_2_21;
output wire [RID_WIDTH-1:0] dout_2_22;
output wire dout_valid_2_22;
output wire [RID_WIDTH-1:0] dout_2_23;
output wire dout_valid_2_23;
output wire [RID_WIDTH-1:0] dout_2_24;
output wire dout_valid_2_24;
output wire [RID_WIDTH-1:0] dout_2_25;
output wire dout_valid_2_25;
output wire [RID_WIDTH-1:0] dout_2_26;
output wire dout_valid_2_26;
output wire [RID_WIDTH-1:0] dout_2_27;
output wire dout_valid_2_27;
output wire [RID_WIDTH-1:0] dout_2_28;
output wire dout_valid_2_28;
output wire [RID_WIDTH-1:0] dout_2_29;
output wire dout_valid_2_29;
output wire [RID_WIDTH-1:0] dout_2_30;
output wire dout_valid_2_30;
output wire [RID_WIDTH-1:0] dout_2_31;
output wire dout_valid_2_31;
output wire [RID_WIDTH-1:0] dout_3_0;
output wire dout_valid_3_0;
output wire [RID_WIDTH-1:0] dout_3_1;
output wire dout_valid_3_1;
output wire [RID_WIDTH-1:0] dout_3_2;
output wire dout_valid_3_2;
output wire [RID_WIDTH-1:0] dout_3_3;
output wire dout_valid_3_3;
output wire [RID_WIDTH-1:0] dout_3_4;
output wire dout_valid_3_4;
output wire [RID_WIDTH-1:0] dout_3_5;
output wire dout_valid_3_5;
output wire [RID_WIDTH-1:0] dout_3_6;
output wire dout_valid_3_6;
output wire [RID_WIDTH-1:0] dout_3_7;
output wire dout_valid_3_7;
output wire [RID_WIDTH-1:0] dout_3_8;
output wire dout_valid_3_8;
output wire [RID_WIDTH-1:0] dout_3_9;
output wire dout_valid_3_9;
output wire [RID_WIDTH-1:0] dout_3_10;
output wire dout_valid_3_10;
output wire [RID_WIDTH-1:0] dout_3_11;
output wire dout_valid_3_11;
output wire [RID_WIDTH-1:0] dout_3_12;
output wire dout_valid_3_12;
output wire [RID_WIDTH-1:0] dout_3_13;
output wire dout_valid_3_13;
output wire [RID_WIDTH-1:0] dout_3_14;
output wire dout_valid_3_14;
output wire [RID_WIDTH-1:0] dout_3_15;
output wire dout_valid_3_15;
output wire [RID_WIDTH-1:0] dout_3_16;
output wire dout_valid_3_16;
output wire [RID_WIDTH-1:0] dout_3_17;
output wire dout_valid_3_17;
output wire [RID_WIDTH-1:0] dout_3_18;
output wire dout_valid_3_18;
output wire [RID_WIDTH-1:0] dout_3_19;
output wire dout_valid_3_19;
output wire [RID_WIDTH-1:0] dout_3_20;
output wire dout_valid_3_20;
output wire [RID_WIDTH-1:0] dout_3_21;
output wire dout_valid_3_21;
output wire [RID_WIDTH-1:0] dout_3_22;
output wire dout_valid_3_22;
output wire [RID_WIDTH-1:0] dout_3_23;
output wire dout_valid_3_23;
output wire [RID_WIDTH-1:0] dout_3_24;
output wire dout_valid_3_24;
output wire [RID_WIDTH-1:0] dout_3_25;
output wire dout_valid_3_25;
output wire [RID_WIDTH-1:0] dout_3_26;
output wire dout_valid_3_26;
output wire [RID_WIDTH-1:0] dout_3_27;
output wire dout_valid_3_27;
output wire [RID_WIDTH-1:0] dout_3_28;
output wire dout_valid_3_28;
output wire [RID_WIDTH-1:0] dout_3_29;
output wire dout_valid_3_29;
output wire [RID_WIDTH-1:0] dout_3_30;
output wire dout_valid_3_30;
output wire [RID_WIDTH-1:0] dout_3_31;
output wire dout_valid_3_31;
output wire [RID_WIDTH-1:0] dout_4_0;
output wire dout_valid_4_0;
output wire [RID_WIDTH-1:0] dout_4_1;
output wire dout_valid_4_1;
output wire [RID_WIDTH-1:0] dout_4_2;
output wire dout_valid_4_2;
output wire [RID_WIDTH-1:0] dout_4_3;
output wire dout_valid_4_3;
output wire [RID_WIDTH-1:0] dout_4_4;
output wire dout_valid_4_4;
output wire [RID_WIDTH-1:0] dout_4_5;
output wire dout_valid_4_5;
output wire [RID_WIDTH-1:0] dout_4_6;
output wire dout_valid_4_6;
output wire [RID_WIDTH-1:0] dout_4_7;
output wire dout_valid_4_7;
output wire [RID_WIDTH-1:0] dout_4_8;
output wire dout_valid_4_8;
output wire [RID_WIDTH-1:0] dout_4_9;
output wire dout_valid_4_9;
output wire [RID_WIDTH-1:0] dout_4_10;
output wire dout_valid_4_10;
output wire [RID_WIDTH-1:0] dout_4_11;
output wire dout_valid_4_11;
output wire [RID_WIDTH-1:0] dout_4_12;
output wire dout_valid_4_12;
output wire [RID_WIDTH-1:0] dout_4_13;
output wire dout_valid_4_13;
output wire [RID_WIDTH-1:0] dout_4_14;
output wire dout_valid_4_14;
output wire [RID_WIDTH-1:0] dout_4_15;
output wire dout_valid_4_15;
output wire [RID_WIDTH-1:0] dout_4_16;
output wire dout_valid_4_16;
output wire [RID_WIDTH-1:0] dout_4_17;
output wire dout_valid_4_17;
output wire [RID_WIDTH-1:0] dout_4_18;
output wire dout_valid_4_18;
output wire [RID_WIDTH-1:0] dout_4_19;
output wire dout_valid_4_19;
output wire [RID_WIDTH-1:0] dout_4_20;
output wire dout_valid_4_20;
output wire [RID_WIDTH-1:0] dout_4_21;
output wire dout_valid_4_21;
output wire [RID_WIDTH-1:0] dout_4_22;
output wire dout_valid_4_22;
output wire [RID_WIDTH-1:0] dout_4_23;
output wire dout_valid_4_23;
output wire [RID_WIDTH-1:0] dout_4_24;
output wire dout_valid_4_24;
output wire [RID_WIDTH-1:0] dout_4_25;
output wire dout_valid_4_25;
output wire [RID_WIDTH-1:0] dout_4_26;
output wire dout_valid_4_26;
output wire [RID_WIDTH-1:0] dout_4_27;
output wire dout_valid_4_27;
output wire [RID_WIDTH-1:0] dout_4_28;
output wire dout_valid_4_28;
output wire [RID_WIDTH-1:0] dout_4_29;
output wire dout_valid_4_29;
output wire [RID_WIDTH-1:0] dout_4_30;
output wire dout_valid_4_30;
output wire [RID_WIDTH-1:0] dout_4_31;
output wire dout_valid_4_31;
output wire [RID_WIDTH-1:0] dout_5_0;
output wire dout_valid_5_0;
output wire [RID_WIDTH-1:0] dout_5_1;
output wire dout_valid_5_1;
output wire [RID_WIDTH-1:0] dout_5_2;
output wire dout_valid_5_2;
output wire [RID_WIDTH-1:0] dout_5_3;
output wire dout_valid_5_3;
output wire [RID_WIDTH-1:0] dout_5_4;
output wire dout_valid_5_4;
output wire [RID_WIDTH-1:0] dout_5_5;
output wire dout_valid_5_5;
output wire [RID_WIDTH-1:0] dout_5_6;
output wire dout_valid_5_6;
output wire [RID_WIDTH-1:0] dout_5_7;
output wire dout_valid_5_7;
output wire [RID_WIDTH-1:0] dout_5_8;
output wire dout_valid_5_8;
output wire [RID_WIDTH-1:0] dout_5_9;
output wire dout_valid_5_9;
output wire [RID_WIDTH-1:0] dout_5_10;
output wire dout_valid_5_10;
output wire [RID_WIDTH-1:0] dout_5_11;
output wire dout_valid_5_11;
output wire [RID_WIDTH-1:0] dout_5_12;
output wire dout_valid_5_12;
output wire [RID_WIDTH-1:0] dout_5_13;
output wire dout_valid_5_13;
output wire [RID_WIDTH-1:0] dout_5_14;
output wire dout_valid_5_14;
output wire [RID_WIDTH-1:0] dout_5_15;
output wire dout_valid_5_15;
output wire [RID_WIDTH-1:0] dout_5_16;
output wire dout_valid_5_16;
output wire [RID_WIDTH-1:0] dout_5_17;
output wire dout_valid_5_17;
output wire [RID_WIDTH-1:0] dout_5_18;
output wire dout_valid_5_18;
output wire [RID_WIDTH-1:0] dout_5_19;
output wire dout_valid_5_19;
output wire [RID_WIDTH-1:0] dout_5_20;
output wire dout_valid_5_20;
output wire [RID_WIDTH-1:0] dout_5_21;
output wire dout_valid_5_21;
output wire [RID_WIDTH-1:0] dout_5_22;
output wire dout_valid_5_22;
output wire [RID_WIDTH-1:0] dout_5_23;
output wire dout_valid_5_23;
output wire [RID_WIDTH-1:0] dout_5_24;
output wire dout_valid_5_24;
output wire [RID_WIDTH-1:0] dout_5_25;
output wire dout_valid_5_25;
output wire [RID_WIDTH-1:0] dout_5_26;
output wire dout_valid_5_26;
output wire [RID_WIDTH-1:0] dout_5_27;
output wire dout_valid_5_27;
output wire [RID_WIDTH-1:0] dout_5_28;
output wire dout_valid_5_28;
output wire [RID_WIDTH-1:0] dout_5_29;
output wire dout_valid_5_29;
output wire [RID_WIDTH-1:0] dout_5_30;
output wire dout_valid_5_30;
output wire [RID_WIDTH-1:0] dout_5_31;
output wire dout_valid_5_31;
output wire [RID_WIDTH-1:0] dout_6_0;
output wire dout_valid_6_0;
output wire [RID_WIDTH-1:0] dout_6_1;
output wire dout_valid_6_1;
output wire [RID_WIDTH-1:0] dout_6_2;
output wire dout_valid_6_2;
output wire [RID_WIDTH-1:0] dout_6_3;
output wire dout_valid_6_3;
output wire [RID_WIDTH-1:0] dout_6_4;
output wire dout_valid_6_4;
output wire [RID_WIDTH-1:0] dout_6_5;
output wire dout_valid_6_5;
output wire [RID_WIDTH-1:0] dout_6_6;
output wire dout_valid_6_6;
output wire [RID_WIDTH-1:0] dout_6_7;
output wire dout_valid_6_7;
output wire [RID_WIDTH-1:0] dout_6_8;
output wire dout_valid_6_8;
output wire [RID_WIDTH-1:0] dout_6_9;
output wire dout_valid_6_9;
output wire [RID_WIDTH-1:0] dout_6_10;
output wire dout_valid_6_10;
output wire [RID_WIDTH-1:0] dout_6_11;
output wire dout_valid_6_11;
output wire [RID_WIDTH-1:0] dout_6_12;
output wire dout_valid_6_12;
output wire [RID_WIDTH-1:0] dout_6_13;
output wire dout_valid_6_13;
output wire [RID_WIDTH-1:0] dout_6_14;
output wire dout_valid_6_14;
output wire [RID_WIDTH-1:0] dout_6_15;
output wire dout_valid_6_15;
output wire [RID_WIDTH-1:0] dout_6_16;
output wire dout_valid_6_16;
output wire [RID_WIDTH-1:0] dout_6_17;
output wire dout_valid_6_17;
output wire [RID_WIDTH-1:0] dout_6_18;
output wire dout_valid_6_18;
output wire [RID_WIDTH-1:0] dout_6_19;
output wire dout_valid_6_19;
output wire [RID_WIDTH-1:0] dout_6_20;
output wire dout_valid_6_20;
output wire [RID_WIDTH-1:0] dout_6_21;
output wire dout_valid_6_21;
output wire [RID_WIDTH-1:0] dout_6_22;
output wire dout_valid_6_22;
output wire [RID_WIDTH-1:0] dout_6_23;
output wire dout_valid_6_23;
output wire [RID_WIDTH-1:0] dout_6_24;
output wire dout_valid_6_24;
output wire [RID_WIDTH-1:0] dout_6_25;
output wire dout_valid_6_25;
output wire [RID_WIDTH-1:0] dout_6_26;
output wire dout_valid_6_26;
output wire [RID_WIDTH-1:0] dout_6_27;
output wire dout_valid_6_27;
output wire [RID_WIDTH-1:0] dout_6_28;
output wire dout_valid_6_28;
output wire [RID_WIDTH-1:0] dout_6_29;
output wire dout_valid_6_29;
output wire [RID_WIDTH-1:0] dout_6_30;
output wire dout_valid_6_30;
output wire [RID_WIDTH-1:0] dout_6_31;
output wire dout_valid_6_31;
output wire [RID_WIDTH-1:0] dout_7_0;
output wire dout_valid_7_0;
output wire [RID_WIDTH-1:0] dout_7_1;
output wire dout_valid_7_1;
output wire [RID_WIDTH-1:0] dout_7_2;
output wire dout_valid_7_2;
output wire [RID_WIDTH-1:0] dout_7_3;
output wire dout_valid_7_3;
output wire [RID_WIDTH-1:0] dout_7_4;
output wire dout_valid_7_4;
output wire [RID_WIDTH-1:0] dout_7_5;
output wire dout_valid_7_5;
output wire [RID_WIDTH-1:0] dout_7_6;
output wire dout_valid_7_6;
output wire [RID_WIDTH-1:0] dout_7_7;
output wire dout_valid_7_7;
output wire [RID_WIDTH-1:0] dout_7_8;
output wire dout_valid_7_8;
output wire [RID_WIDTH-1:0] dout_7_9;
output wire dout_valid_7_9;
output wire [RID_WIDTH-1:0] dout_7_10;
output wire dout_valid_7_10;
output wire [RID_WIDTH-1:0] dout_7_11;
output wire dout_valid_7_11;
output wire [RID_WIDTH-1:0] dout_7_12;
output wire dout_valid_7_12;
output wire [RID_WIDTH-1:0] dout_7_13;
output wire dout_valid_7_13;
output wire [RID_WIDTH-1:0] dout_7_14;
output wire dout_valid_7_14;
output wire [RID_WIDTH-1:0] dout_7_15;
output wire dout_valid_7_15;
output wire [RID_WIDTH-1:0] dout_7_16;
output wire dout_valid_7_16;
output wire [RID_WIDTH-1:0] dout_7_17;
output wire dout_valid_7_17;
output wire [RID_WIDTH-1:0] dout_7_18;
output wire dout_valid_7_18;
output wire [RID_WIDTH-1:0] dout_7_19;
output wire dout_valid_7_19;
output wire [RID_WIDTH-1:0] dout_7_20;
output wire dout_valid_7_20;
output wire [RID_WIDTH-1:0] dout_7_21;
output wire dout_valid_7_21;
output wire [RID_WIDTH-1:0] dout_7_22;
output wire dout_valid_7_22;
output wire [RID_WIDTH-1:0] dout_7_23;
output wire dout_valid_7_23;
output wire [RID_WIDTH-1:0] dout_7_24;
output wire dout_valid_7_24;
output wire [RID_WIDTH-1:0] dout_7_25;
output wire dout_valid_7_25;
output wire [RID_WIDTH-1:0] dout_7_26;
output wire dout_valid_7_26;
output wire [RID_WIDTH-1:0] dout_7_27;
output wire dout_valid_7_27;
output wire [RID_WIDTH-1:0] dout_7_28;
output wire dout_valid_7_28;
output wire [RID_WIDTH-1:0] dout_7_29;
output wire dout_valid_7_29;
output wire [RID_WIDTH-1:0] dout_7_30;
output wire dout_valid_7_30;
output wire [RID_WIDTH-1:0] dout_7_31;
output wire dout_valid_7_31;

reg  [15-1:0] addr_0_0;
wire din_valid_0_0;
wire addr_valid_0_0;
reg  [15-1:0] addr_0_1;
wire din_valid_0_1;
wire addr_valid_0_1;
reg  [15-1:0] addr_0_2;
wire din_valid_0_2;
wire addr_valid_0_2;
reg  [15-1:0] addr_0_3;
wire din_valid_0_3;
wire addr_valid_0_3;
reg  [15-1:0] addr_0_4;
wire din_valid_0_4;
wire addr_valid_0_4;
reg  [15-1:0] addr_0_5;
wire din_valid_0_5;
wire addr_valid_0_5;
reg  [15-1:0] addr_0_6;
wire din_valid_0_6;
wire addr_valid_0_6;
reg  [15-1:0] addr_0_7;
wire din_valid_0_7;
wire addr_valid_0_7;
reg  [15-1:0] addr_0_8;
wire din_valid_0_8;
wire addr_valid_0_8;
reg  [15-1:0] addr_0_9;
wire din_valid_0_9;
wire addr_valid_0_9;
reg  [15-1:0] addr_0_10;
wire din_valid_0_10;
wire addr_valid_0_10;
reg  [15-1:0] addr_0_11;
wire din_valid_0_11;
wire addr_valid_0_11;
reg  [15-1:0] addr_0_12;
wire din_valid_0_12;
wire addr_valid_0_12;
reg  [15-1:0] addr_0_13;
wire din_valid_0_13;
wire addr_valid_0_13;
reg  [15-1:0] addr_0_14;
wire din_valid_0_14;
wire addr_valid_0_14;
reg  [15-1:0] addr_0_15;
wire din_valid_0_15;
wire addr_valid_0_15;
reg  [15-1:0] addr_0_16;
wire din_valid_0_16;
wire addr_valid_0_16;
reg  [15-1:0] addr_0_17;
wire din_valid_0_17;
wire addr_valid_0_17;
reg  [15-1:0] addr_0_18;
wire din_valid_0_18;
wire addr_valid_0_18;
reg  [15-1:0] addr_0_19;
wire din_valid_0_19;
wire addr_valid_0_19;
reg  [15-1:0] addr_0_20;
wire din_valid_0_20;
wire addr_valid_0_20;
reg  [15-1:0] addr_0_21;
wire din_valid_0_21;
wire addr_valid_0_21;
reg  [15-1:0] addr_0_22;
wire din_valid_0_22;
wire addr_valid_0_22;
reg  [15-1:0] addr_0_23;
wire din_valid_0_23;
wire addr_valid_0_23;
reg  [15-1:0] addr_0_24;
wire din_valid_0_24;
wire addr_valid_0_24;
reg  [15-1:0] addr_0_25;
wire din_valid_0_25;
wire addr_valid_0_25;
reg  [15-1:0] addr_0_26;
wire din_valid_0_26;
wire addr_valid_0_26;
reg  [15-1:0] addr_0_27;
wire din_valid_0_27;
wire addr_valid_0_27;
reg  [15-1:0] addr_0_28;
wire din_valid_0_28;
wire addr_valid_0_28;
reg  [15-1:0] addr_0_29;
wire din_valid_0_29;
wire addr_valid_0_29;
reg  [15-1:0] addr_0_30;
wire din_valid_0_30;
wire addr_valid_0_30;
reg  [15-1:0] addr_0_31;
wire din_valid_0_31;
wire addr_valid_0_31;
reg  [15-1:0] addr_1_0;
wire din_valid_1_0;
wire addr_valid_1_0;
reg  [15-1:0] addr_1_1;
wire din_valid_1_1;
wire addr_valid_1_1;
reg  [15-1:0] addr_1_2;
wire din_valid_1_2;
wire addr_valid_1_2;
reg  [15-1:0] addr_1_3;
wire din_valid_1_3;
wire addr_valid_1_3;
reg  [15-1:0] addr_1_4;
wire din_valid_1_4;
wire addr_valid_1_4;
reg  [15-1:0] addr_1_5;
wire din_valid_1_5;
wire addr_valid_1_5;
reg  [15-1:0] addr_1_6;
wire din_valid_1_6;
wire addr_valid_1_6;
reg  [15-1:0] addr_1_7;
wire din_valid_1_7;
wire addr_valid_1_7;
reg  [15-1:0] addr_1_8;
wire din_valid_1_8;
wire addr_valid_1_8;
reg  [15-1:0] addr_1_9;
wire din_valid_1_9;
wire addr_valid_1_9;
reg  [15-1:0] addr_1_10;
wire din_valid_1_10;
wire addr_valid_1_10;
reg  [15-1:0] addr_1_11;
wire din_valid_1_11;
wire addr_valid_1_11;
reg  [15-1:0] addr_1_12;
wire din_valid_1_12;
wire addr_valid_1_12;
reg  [15-1:0] addr_1_13;
wire din_valid_1_13;
wire addr_valid_1_13;
reg  [15-1:0] addr_1_14;
wire din_valid_1_14;
wire addr_valid_1_14;
reg  [15-1:0] addr_1_15;
wire din_valid_1_15;
wire addr_valid_1_15;
reg  [15-1:0] addr_1_16;
wire din_valid_1_16;
wire addr_valid_1_16;
reg  [15-1:0] addr_1_17;
wire din_valid_1_17;
wire addr_valid_1_17;
reg  [15-1:0] addr_1_18;
wire din_valid_1_18;
wire addr_valid_1_18;
reg  [15-1:0] addr_1_19;
wire din_valid_1_19;
wire addr_valid_1_19;
reg  [15-1:0] addr_1_20;
wire din_valid_1_20;
wire addr_valid_1_20;
reg  [15-1:0] addr_1_21;
wire din_valid_1_21;
wire addr_valid_1_21;
reg  [15-1:0] addr_1_22;
wire din_valid_1_22;
wire addr_valid_1_22;
reg  [15-1:0] addr_1_23;
wire din_valid_1_23;
wire addr_valid_1_23;
reg  [15-1:0] addr_1_24;
wire din_valid_1_24;
wire addr_valid_1_24;
reg  [15-1:0] addr_1_25;
wire din_valid_1_25;
wire addr_valid_1_25;
reg  [15-1:0] addr_1_26;
wire din_valid_1_26;
wire addr_valid_1_26;
reg  [15-1:0] addr_1_27;
wire din_valid_1_27;
wire addr_valid_1_27;
reg  [15-1:0] addr_1_28;
wire din_valid_1_28;
wire addr_valid_1_28;
reg  [15-1:0] addr_1_29;
wire din_valid_1_29;
wire addr_valid_1_29;
reg  [15-1:0] addr_1_30;
wire din_valid_1_30;
wire addr_valid_1_30;
reg  [15-1:0] addr_1_31;
wire din_valid_1_31;
wire addr_valid_1_31;
reg  [12-1:0] addr_2_0;
wire din_valid_2_0;
wire addr_valid_2_0;
reg  [12-1:0] addr_2_1;
wire din_valid_2_1;
wire addr_valid_2_1;
reg  [12-1:0] addr_2_2;
wire din_valid_2_2;
wire addr_valid_2_2;
reg  [12-1:0] addr_2_3;
wire din_valid_2_3;
wire addr_valid_2_3;
reg  [12-1:0] addr_2_4;
wire din_valid_2_4;
wire addr_valid_2_4;
reg  [12-1:0] addr_2_5;
wire din_valid_2_5;
wire addr_valid_2_5;
reg  [12-1:0] addr_2_6;
wire din_valid_2_6;
wire addr_valid_2_6;
reg  [12-1:0] addr_2_7;
wire din_valid_2_7;
wire addr_valid_2_7;
reg  [12-1:0] addr_2_8;
wire din_valid_2_8;
wire addr_valid_2_8;
reg  [12-1:0] addr_2_9;
wire din_valid_2_9;
wire addr_valid_2_9;
reg  [12-1:0] addr_2_10;
wire din_valid_2_10;
wire addr_valid_2_10;
reg  [12-1:0] addr_2_11;
wire din_valid_2_11;
wire addr_valid_2_11;
reg  [12-1:0] addr_2_12;
wire din_valid_2_12;
wire addr_valid_2_12;
reg  [12-1:0] addr_2_13;
wire din_valid_2_13;
wire addr_valid_2_13;
reg  [12-1:0] addr_2_14;
wire din_valid_2_14;
wire addr_valid_2_14;
reg  [12-1:0] addr_2_15;
wire din_valid_2_15;
wire addr_valid_2_15;
reg  [12-1:0] addr_2_16;
wire din_valid_2_16;
wire addr_valid_2_16;
reg  [12-1:0] addr_2_17;
wire din_valid_2_17;
wire addr_valid_2_17;
reg  [12-1:0] addr_2_18;
wire din_valid_2_18;
wire addr_valid_2_18;
reg  [12-1:0] addr_2_19;
wire din_valid_2_19;
wire addr_valid_2_19;
reg  [12-1:0] addr_2_20;
wire din_valid_2_20;
wire addr_valid_2_20;
reg  [12-1:0] addr_2_21;
wire din_valid_2_21;
wire addr_valid_2_21;
reg  [12-1:0] addr_2_22;
wire din_valid_2_22;
wire addr_valid_2_22;
reg  [12-1:0] addr_2_23;
wire din_valid_2_23;
wire addr_valid_2_23;
reg  [12-1:0] addr_2_24;
wire din_valid_2_24;
wire addr_valid_2_24;
reg  [12-1:0] addr_2_25;
wire din_valid_2_25;
wire addr_valid_2_25;
reg  [12-1:0] addr_2_26;
wire din_valid_2_26;
wire addr_valid_2_26;
reg  [12-1:0] addr_2_27;
wire din_valid_2_27;
wire addr_valid_2_27;
reg  [12-1:0] addr_2_28;
wire din_valid_2_28;
wire addr_valid_2_28;
reg  [12-1:0] addr_2_29;
wire din_valid_2_29;
wire addr_valid_2_29;
reg  [12-1:0] addr_2_30;
wire din_valid_2_30;
wire addr_valid_2_30;
reg  [12-1:0] addr_2_31;
wire din_valid_2_31;
wire addr_valid_2_31;
reg  [12-1:0] addr_3_0;
wire din_valid_3_0;
wire addr_valid_3_0;
reg  [12-1:0] addr_3_1;
wire din_valid_3_1;
wire addr_valid_3_1;
reg  [12-1:0] addr_3_2;
wire din_valid_3_2;
wire addr_valid_3_2;
reg  [12-1:0] addr_3_3;
wire din_valid_3_3;
wire addr_valid_3_3;
reg  [12-1:0] addr_3_4;
wire din_valid_3_4;
wire addr_valid_3_4;
reg  [12-1:0] addr_3_5;
wire din_valid_3_5;
wire addr_valid_3_5;
reg  [12-1:0] addr_3_6;
wire din_valid_3_6;
wire addr_valid_3_6;
reg  [12-1:0] addr_3_7;
wire din_valid_3_7;
wire addr_valid_3_7;
reg  [12-1:0] addr_3_8;
wire din_valid_3_8;
wire addr_valid_3_8;
reg  [12-1:0] addr_3_9;
wire din_valid_3_9;
wire addr_valid_3_9;
reg  [12-1:0] addr_3_10;
wire din_valid_3_10;
wire addr_valid_3_10;
reg  [12-1:0] addr_3_11;
wire din_valid_3_11;
wire addr_valid_3_11;
reg  [12-1:0] addr_3_12;
wire din_valid_3_12;
wire addr_valid_3_12;
reg  [12-1:0] addr_3_13;
wire din_valid_3_13;
wire addr_valid_3_13;
reg  [12-1:0] addr_3_14;
wire din_valid_3_14;
wire addr_valid_3_14;
reg  [12-1:0] addr_3_15;
wire din_valid_3_15;
wire addr_valid_3_15;
reg  [12-1:0] addr_3_16;
wire din_valid_3_16;
wire addr_valid_3_16;
reg  [12-1:0] addr_3_17;
wire din_valid_3_17;
wire addr_valid_3_17;
reg  [12-1:0] addr_3_18;
wire din_valid_3_18;
wire addr_valid_3_18;
reg  [12-1:0] addr_3_19;
wire din_valid_3_19;
wire addr_valid_3_19;
reg  [12-1:0] addr_3_20;
wire din_valid_3_20;
wire addr_valid_3_20;
reg  [12-1:0] addr_3_21;
wire din_valid_3_21;
wire addr_valid_3_21;
reg  [12-1:0] addr_3_22;
wire din_valid_3_22;
wire addr_valid_3_22;
reg  [12-1:0] addr_3_23;
wire din_valid_3_23;
wire addr_valid_3_23;
reg  [12-1:0] addr_3_24;
wire din_valid_3_24;
wire addr_valid_3_24;
reg  [12-1:0] addr_3_25;
wire din_valid_3_25;
wire addr_valid_3_25;
reg  [12-1:0] addr_3_26;
wire din_valid_3_26;
wire addr_valid_3_26;
reg  [12-1:0] addr_3_27;
wire din_valid_3_27;
wire addr_valid_3_27;
reg  [12-1:0] addr_3_28;
wire din_valid_3_28;
wire addr_valid_3_28;
reg  [12-1:0] addr_3_29;
wire din_valid_3_29;
wire addr_valid_3_29;
reg  [12-1:0] addr_3_30;
wire din_valid_3_30;
wire addr_valid_3_30;
reg  [12-1:0] addr_3_31;
wire din_valid_3_31;
wire addr_valid_3_31;
reg  [11-1:0] addr_4_0;
wire din_valid_4_0;
wire addr_valid_4_0;
reg  [11-1:0] addr_4_1;
wire din_valid_4_1;
wire addr_valid_4_1;
reg  [11-1:0] addr_4_2;
wire din_valid_4_2;
wire addr_valid_4_2;
reg  [11-1:0] addr_4_3;
wire din_valid_4_3;
wire addr_valid_4_3;
reg  [11-1:0] addr_4_4;
wire din_valid_4_4;
wire addr_valid_4_4;
reg  [11-1:0] addr_4_5;
wire din_valid_4_5;
wire addr_valid_4_5;
reg  [11-1:0] addr_4_6;
wire din_valid_4_6;
wire addr_valid_4_6;
reg  [11-1:0] addr_4_7;
wire din_valid_4_7;
wire addr_valid_4_7;
reg  [11-1:0] addr_4_8;
wire din_valid_4_8;
wire addr_valid_4_8;
reg  [11-1:0] addr_4_9;
wire din_valid_4_9;
wire addr_valid_4_9;
reg  [11-1:0] addr_4_10;
wire din_valid_4_10;
wire addr_valid_4_10;
reg  [11-1:0] addr_4_11;
wire din_valid_4_11;
wire addr_valid_4_11;
reg  [11-1:0] addr_4_12;
wire din_valid_4_12;
wire addr_valid_4_12;
reg  [11-1:0] addr_4_13;
wire din_valid_4_13;
wire addr_valid_4_13;
reg  [11-1:0] addr_4_14;
wire din_valid_4_14;
wire addr_valid_4_14;
reg  [11-1:0] addr_4_15;
wire din_valid_4_15;
wire addr_valid_4_15;
reg  [11-1:0] addr_4_16;
wire din_valid_4_16;
wire addr_valid_4_16;
reg  [11-1:0] addr_4_17;
wire din_valid_4_17;
wire addr_valid_4_17;
reg  [11-1:0] addr_4_18;
wire din_valid_4_18;
wire addr_valid_4_18;
reg  [11-1:0] addr_4_19;
wire din_valid_4_19;
wire addr_valid_4_19;
reg  [11-1:0] addr_4_20;
wire din_valid_4_20;
wire addr_valid_4_20;
reg  [11-1:0] addr_4_21;
wire din_valid_4_21;
wire addr_valid_4_21;
reg  [11-1:0] addr_4_22;
wire din_valid_4_22;
wire addr_valid_4_22;
reg  [11-1:0] addr_4_23;
wire din_valid_4_23;
wire addr_valid_4_23;
reg  [11-1:0] addr_4_24;
wire din_valid_4_24;
wire addr_valid_4_24;
reg  [11-1:0] addr_4_25;
wire din_valid_4_25;
wire addr_valid_4_25;
reg  [11-1:0] addr_4_26;
wire din_valid_4_26;
wire addr_valid_4_26;
reg  [11-1:0] addr_4_27;
wire din_valid_4_27;
wire addr_valid_4_27;
reg  [11-1:0] addr_4_28;
wire din_valid_4_28;
wire addr_valid_4_28;
reg  [11-1:0] addr_4_29;
wire din_valid_4_29;
wire addr_valid_4_29;
reg  [11-1:0] addr_4_30;
wire din_valid_4_30;
wire addr_valid_4_30;
reg  [11-1:0] addr_4_31;
wire din_valid_4_31;
wire addr_valid_4_31;
reg  [12-1:0] addr_5_0;
wire din_valid_5_0;
wire addr_valid_5_0;
reg  [12-1:0] addr_5_1;
wire din_valid_5_1;
wire addr_valid_5_1;
reg  [12-1:0] addr_5_2;
wire din_valid_5_2;
wire addr_valid_5_2;
reg  [12-1:0] addr_5_3;
wire din_valid_5_3;
wire addr_valid_5_3;
reg  [12-1:0] addr_5_4;
wire din_valid_5_4;
wire addr_valid_5_4;
reg  [12-1:0] addr_5_5;
wire din_valid_5_5;
wire addr_valid_5_5;
reg  [12-1:0] addr_5_6;
wire din_valid_5_6;
wire addr_valid_5_6;
reg  [12-1:0] addr_5_7;
wire din_valid_5_7;
wire addr_valid_5_7;
reg  [12-1:0] addr_5_8;
wire din_valid_5_8;
wire addr_valid_5_8;
reg  [12-1:0] addr_5_9;
wire din_valid_5_9;
wire addr_valid_5_9;
reg  [12-1:0] addr_5_10;
wire din_valid_5_10;
wire addr_valid_5_10;
reg  [12-1:0] addr_5_11;
wire din_valid_5_11;
wire addr_valid_5_11;
reg  [12-1:0] addr_5_12;
wire din_valid_5_12;
wire addr_valid_5_12;
reg  [12-1:0] addr_5_13;
wire din_valid_5_13;
wire addr_valid_5_13;
reg  [12-1:0] addr_5_14;
wire din_valid_5_14;
wire addr_valid_5_14;
reg  [12-1:0] addr_5_15;
wire din_valid_5_15;
wire addr_valid_5_15;
reg  [12-1:0] addr_5_16;
wire din_valid_5_16;
wire addr_valid_5_16;
reg  [12-1:0] addr_5_17;
wire din_valid_5_17;
wire addr_valid_5_17;
reg  [12-1:0] addr_5_18;
wire din_valid_5_18;
wire addr_valid_5_18;
reg  [12-1:0] addr_5_19;
wire din_valid_5_19;
wire addr_valid_5_19;
reg  [12-1:0] addr_5_20;
wire din_valid_5_20;
wire addr_valid_5_20;
reg  [12-1:0] addr_5_21;
wire din_valid_5_21;
wire addr_valid_5_21;
reg  [12-1:0] addr_5_22;
wire din_valid_5_22;
wire addr_valid_5_22;
reg  [12-1:0] addr_5_23;
wire din_valid_5_23;
wire addr_valid_5_23;
reg  [12-1:0] addr_5_24;
wire din_valid_5_24;
wire addr_valid_5_24;
reg  [12-1:0] addr_5_25;
wire din_valid_5_25;
wire addr_valid_5_25;
reg  [12-1:0] addr_5_26;
wire din_valid_5_26;
wire addr_valid_5_26;
reg  [12-1:0] addr_5_27;
wire din_valid_5_27;
wire addr_valid_5_27;
reg  [12-1:0] addr_5_28;
wire din_valid_5_28;
wire addr_valid_5_28;
reg  [12-1:0] addr_5_29;
wire din_valid_5_29;
wire addr_valid_5_29;
reg  [12-1:0] addr_5_30;
wire din_valid_5_30;
wire addr_valid_5_30;
reg  [12-1:0] addr_5_31;
wire din_valid_5_31;
wire addr_valid_5_31;
reg  [10-1:0] addr_6_0;
wire din_valid_6_0;
wire addr_valid_6_0;
reg  [10-1:0] addr_6_1;
wire din_valid_6_1;
wire addr_valid_6_1;
reg  [10-1:0] addr_6_2;
wire din_valid_6_2;
wire addr_valid_6_2;
reg  [10-1:0] addr_6_3;
wire din_valid_6_3;
wire addr_valid_6_3;
reg  [10-1:0] addr_6_4;
wire din_valid_6_4;
wire addr_valid_6_4;
reg  [10-1:0] addr_6_5;
wire din_valid_6_5;
wire addr_valid_6_5;
reg  [10-1:0] addr_6_6;
wire din_valid_6_6;
wire addr_valid_6_6;
reg  [10-1:0] addr_6_7;
wire din_valid_6_7;
wire addr_valid_6_7;
reg  [10-1:0] addr_6_8;
wire din_valid_6_8;
wire addr_valid_6_8;
reg  [10-1:0] addr_6_9;
wire din_valid_6_9;
wire addr_valid_6_9;
reg  [10-1:0] addr_6_10;
wire din_valid_6_10;
wire addr_valid_6_10;
reg  [10-1:0] addr_6_11;
wire din_valid_6_11;
wire addr_valid_6_11;
reg  [10-1:0] addr_6_12;
wire din_valid_6_12;
wire addr_valid_6_12;
reg  [10-1:0] addr_6_13;
wire din_valid_6_13;
wire addr_valid_6_13;
reg  [10-1:0] addr_6_14;
wire din_valid_6_14;
wire addr_valid_6_14;
reg  [10-1:0] addr_6_15;
wire din_valid_6_15;
wire addr_valid_6_15;
reg  [10-1:0] addr_6_16;
wire din_valid_6_16;
wire addr_valid_6_16;
reg  [10-1:0] addr_6_17;
wire din_valid_6_17;
wire addr_valid_6_17;
reg  [10-1:0] addr_6_18;
wire din_valid_6_18;
wire addr_valid_6_18;
reg  [10-1:0] addr_6_19;
wire din_valid_6_19;
wire addr_valid_6_19;
reg  [10-1:0] addr_6_20;
wire din_valid_6_20;
wire addr_valid_6_20;
reg  [10-1:0] addr_6_21;
wire din_valid_6_21;
wire addr_valid_6_21;
reg  [10-1:0] addr_6_22;
wire din_valid_6_22;
wire addr_valid_6_22;
reg  [10-1:0] addr_6_23;
wire din_valid_6_23;
wire addr_valid_6_23;
reg  [10-1:0] addr_6_24;
wire din_valid_6_24;
wire addr_valid_6_24;
reg  [10-1:0] addr_6_25;
wire din_valid_6_25;
wire addr_valid_6_25;
reg  [10-1:0] addr_6_26;
wire din_valid_6_26;
wire addr_valid_6_26;
reg  [10-1:0] addr_6_27;
wire din_valid_6_27;
wire addr_valid_6_27;
reg  [10-1:0] addr_6_28;
wire din_valid_6_28;
wire addr_valid_6_28;
reg  [10-1:0] addr_6_29;
wire din_valid_6_29;
wire addr_valid_6_29;
reg  [10-1:0] addr_6_30;
wire din_valid_6_30;
wire addr_valid_6_30;
reg  [10-1:0] addr_6_31;
wire din_valid_6_31;
wire addr_valid_6_31;
reg  [8-1:0] addr_7_0;
wire din_valid_7_0;
wire addr_valid_7_0;
reg  [8-1:0] addr_7_1;
wire din_valid_7_1;
wire addr_valid_7_1;
reg  [8-1:0] addr_7_2;
wire din_valid_7_2;
wire addr_valid_7_2;
reg  [8-1:0] addr_7_3;
wire din_valid_7_3;
wire addr_valid_7_3;
reg  [8-1:0] addr_7_4;
wire din_valid_7_4;
wire addr_valid_7_4;
reg  [8-1:0] addr_7_5;
wire din_valid_7_5;
wire addr_valid_7_5;
reg  [8-1:0] addr_7_6;
wire din_valid_7_6;
wire addr_valid_7_6;
reg  [8-1:0] addr_7_7;
wire din_valid_7_7;
wire addr_valid_7_7;
reg  [8-1:0] addr_7_8;
wire din_valid_7_8;
wire addr_valid_7_8;
reg  [8-1:0] addr_7_9;
wire din_valid_7_9;
wire addr_valid_7_9;
reg  [8-1:0] addr_7_10;
wire din_valid_7_10;
wire addr_valid_7_10;
reg  [8-1:0] addr_7_11;
wire din_valid_7_11;
wire addr_valid_7_11;
reg  [8-1:0] addr_7_12;
wire din_valid_7_12;
wire addr_valid_7_12;
reg  [8-1:0] addr_7_13;
wire din_valid_7_13;
wire addr_valid_7_13;
reg  [8-1:0] addr_7_14;
wire din_valid_7_14;
wire addr_valid_7_14;
reg  [8-1:0] addr_7_15;
wire din_valid_7_15;
wire addr_valid_7_15;
reg  [8-1:0] addr_7_16;
wire din_valid_7_16;
wire addr_valid_7_16;
reg  [8-1:0] addr_7_17;
wire din_valid_7_17;
wire addr_valid_7_17;
reg  [8-1:0] addr_7_18;
wire din_valid_7_18;
wire addr_valid_7_18;
reg  [8-1:0] addr_7_19;
wire din_valid_7_19;
wire addr_valid_7_19;
reg  [8-1:0] addr_7_20;
wire din_valid_7_20;
wire addr_valid_7_20;
reg  [8-1:0] addr_7_21;
wire din_valid_7_21;
wire addr_valid_7_21;
reg  [8-1:0] addr_7_22;
wire din_valid_7_22;
wire addr_valid_7_22;
reg  [8-1:0] addr_7_23;
wire din_valid_7_23;
wire addr_valid_7_23;
reg  [8-1:0] addr_7_24;
wire din_valid_7_24;
wire addr_valid_7_24;
reg  [8-1:0] addr_7_25;
wire din_valid_7_25;
wire addr_valid_7_25;
reg  [8-1:0] addr_7_26;
wire din_valid_7_26;
wire addr_valid_7_26;
reg  [8-1:0] addr_7_27;
wire din_valid_7_27;
wire addr_valid_7_27;
reg  [8-1:0] addr_7_28;
wire din_valid_7_28;
wire addr_valid_7_28;
reg  [8-1:0] addr_7_29;
wire din_valid_7_29;
wire addr_valid_7_29;
reg  [8-1:0] addr_7_30;
wire din_valid_7_30;
wire addr_valid_7_30;
reg  [8-1:0] addr_7_31;
wire din_valid_7_31;
wire addr_valid_7_31;

reg [63:0] din_reg;
reg din_valid_reg;

// Doing all necessary multiplies per double_byte
wire [(32+7)*8-1:0] padded_din;
wire [32-1:0] din_signs;
wire [32-1:0] din_signs_reg;

wire [31:0] din_0_ab0;
wire [31:0] din_0_ab1;
wire [31:0] din_0_ab2;
wire [31:0] din_0_ab3;
wire [31:0] din_0_ab0_1sc;
wire [31:0] din_0_ab1_1sc;
wire [31:0] din_0_ab2_1sc;
wire [31:0] din_0_ab3_1sc;
wire [23:0] din_0_msk_ab0;
wire [23:0] din_0_msk_ab1;
wire [23:0] din_0_msk_ab2;
wire [23:0] din_0_msk_ab3;
wire [23:0] din_0_msk_ab0_1sc;
wire [23:0] din_0_msk_ab1_1sc;
wire [23:0] din_0_msk_ab2_1sc;
wire [23:0] din_0_msk_ab3_1sc;
wire [31:0] din_1_ab0;
wire [31:0] din_1_ab1;
wire [31:0] din_1_ab2;
wire [31:0] din_1_ab3;
wire [31:0] din_1_ab0_1sc;
wire [31:0] din_1_ab1_1sc;
wire [31:0] din_1_ab2_1sc;
wire [31:0] din_1_ab3_1sc;
wire [23:0] din_1_msk_ab0;
wire [23:0] din_1_msk_ab1;
wire [23:0] din_1_msk_ab2;
wire [23:0] din_1_msk_ab3;
wire [23:0] din_1_msk_ab0_1sc;
wire [23:0] din_1_msk_ab1_1sc;
wire [23:0] din_1_msk_ab2_1sc;
wire [23:0] din_1_msk_ab3_1sc;
wire [31:0] din_2_ab0;
wire [31:0] din_2_ab1;
wire [31:0] din_2_ab2;
wire [31:0] din_2_ab3;
wire [31:0] din_2_ab0_1sc;
wire [31:0] din_2_ab1_1sc;
wire [31:0] din_2_ab2_1sc;
wire [31:0] din_2_ab3_1sc;
wire [23:0] din_2_msk_ab0;
wire [23:0] din_2_msk_ab1;
wire [23:0] din_2_msk_ab2;
wire [23:0] din_2_msk_ab3;
wire [23:0] din_2_msk_ab0_1sc;
wire [23:0] din_2_msk_ab1_1sc;
wire [23:0] din_2_msk_ab2_1sc;
wire [23:0] din_2_msk_ab3_1sc;
wire [31:0] din_3_ab0;
wire [31:0] din_3_ab1;
wire [31:0] din_3_ab2;
wire [31:0] din_3_ab3;
wire [31:0] din_3_ab0_1sc;
wire [31:0] din_3_ab1_1sc;
wire [31:0] din_3_ab2_1sc;
wire [31:0] din_3_ab3_1sc;
wire [23:0] din_3_msk_ab0;
wire [23:0] din_3_msk_ab1;
wire [23:0] din_3_msk_ab2;
wire [23:0] din_3_msk_ab3;
wire [23:0] din_3_msk_ab0_1sc;
wire [23:0] din_3_msk_ab1_1sc;
wire [23:0] din_3_msk_ab2_1sc;
wire [23:0] din_3_msk_ab3_1sc;
wire [31:0] din_4_ab0;
wire [31:0] din_4_ab1;
wire [31:0] din_4_ab2;
wire [31:0] din_4_ab3;
wire [31:0] din_4_ab0_1sc;
wire [31:0] din_4_ab1_1sc;
wire [31:0] din_4_ab2_1sc;
wire [31:0] din_4_ab3_1sc;
wire [23:0] din_4_msk_ab0;
wire [23:0] din_4_msk_ab1;
wire [23:0] din_4_msk_ab2;
wire [23:0] din_4_msk_ab3;
wire [23:0] din_4_msk_ab0_1sc;
wire [23:0] din_4_msk_ab1_1sc;
wire [23:0] din_4_msk_ab2_1sc;
wire [23:0] din_4_msk_ab3_1sc;
wire [31:0] din_5_ab0;
wire [31:0] din_5_ab1;
wire [31:0] din_5_ab2;
wire [31:0] din_5_ab3;
wire [31:0] din_5_ab0_1sc;
wire [31:0] din_5_ab1_1sc;
wire [31:0] din_5_ab2_1sc;
wire [31:0] din_5_ab3_1sc;
wire [23:0] din_5_msk_ab0;
wire [23:0] din_5_msk_ab1;
wire [23:0] din_5_msk_ab2;
wire [23:0] din_5_msk_ab3;
wire [23:0] din_5_msk_ab0_1sc;
wire [23:0] din_5_msk_ab1_1sc;
wire [23:0] din_5_msk_ab2_1sc;
wire [23:0] din_5_msk_ab3_1sc;
wire [31:0] din_6_ab0;
wire [31:0] din_6_ab1;
wire [31:0] din_6_ab2;
wire [31:0] din_6_ab3;
wire [31:0] din_6_ab0_1sc;
wire [31:0] din_6_ab1_1sc;
wire [31:0] din_6_ab2_1sc;
wire [31:0] din_6_ab3_1sc;
wire [23:0] din_6_msk_ab0;
wire [23:0] din_6_msk_ab1;
wire [23:0] din_6_msk_ab2;
wire [23:0] din_6_msk_ab3;
wire [23:0] din_6_msk_ab0_1sc;
wire [23:0] din_6_msk_ab1_1sc;
wire [23:0] din_6_msk_ab2_1sc;
wire [23:0] din_6_msk_ab3_1sc;
wire [31:0] din_7_ab0;
wire [31:0] din_7_ab1;
wire [31:0] din_7_ab2;
wire [31:0] din_7_ab3;
wire [31:0] din_7_ab0_1sc;
wire [31:0] din_7_ab1_1sc;
wire [31:0] din_7_ab2_1sc;
wire [31:0] din_7_ab3_1sc;
wire [23:0] din_7_msk_ab0;
wire [23:0] din_7_msk_ab1;
wire [23:0] din_7_msk_ab2;
wire [23:0] din_7_msk_ab3;
wire [23:0] din_7_msk_ab0_1sc;
wire [23:0] din_7_msk_ab1_1sc;
wire [23:0] din_7_msk_ab2_1sc;
wire [23:0] din_7_msk_ab3_1sc;
wire [31:0] din_8_ab0;
wire [31:0] din_8_ab1;
wire [31:0] din_8_ab2;
wire [31:0] din_8_ab3;
wire [31:0] din_8_ab0_1sc;
wire [31:0] din_8_ab1_1sc;
wire [31:0] din_8_ab2_1sc;
wire [31:0] din_8_ab3_1sc;
wire [23:0] din_8_msk_ab0;
wire [23:0] din_8_msk_ab1;
wire [23:0] din_8_msk_ab2;
wire [23:0] din_8_msk_ab3;
wire [23:0] din_8_msk_ab0_1sc;
wire [23:0] din_8_msk_ab1_1sc;
wire [23:0] din_8_msk_ab2_1sc;
wire [23:0] din_8_msk_ab3_1sc;
wire [31:0] din_9_ab0;
wire [31:0] din_9_ab1;
wire [31:0] din_9_ab2;
wire [31:0] din_9_ab3;
wire [31:0] din_9_ab0_1sc;
wire [31:0] din_9_ab1_1sc;
wire [31:0] din_9_ab2_1sc;
wire [31:0] din_9_ab3_1sc;
wire [23:0] din_9_msk_ab0;
wire [23:0] din_9_msk_ab1;
wire [23:0] din_9_msk_ab2;
wire [23:0] din_9_msk_ab3;
wire [23:0] din_9_msk_ab0_1sc;
wire [23:0] din_9_msk_ab1_1sc;
wire [23:0] din_9_msk_ab2_1sc;
wire [23:0] din_9_msk_ab3_1sc;
wire [31:0] din_10_ab0;
wire [31:0] din_10_ab1;
wire [31:0] din_10_ab2;
wire [31:0] din_10_ab3;
wire [31:0] din_10_ab0_1sc;
wire [31:0] din_10_ab1_1sc;
wire [31:0] din_10_ab2_1sc;
wire [31:0] din_10_ab3_1sc;
wire [23:0] din_10_msk_ab0;
wire [23:0] din_10_msk_ab1;
wire [23:0] din_10_msk_ab2;
wire [23:0] din_10_msk_ab3;
wire [23:0] din_10_msk_ab0_1sc;
wire [23:0] din_10_msk_ab1_1sc;
wire [23:0] din_10_msk_ab2_1sc;
wire [23:0] din_10_msk_ab3_1sc;
wire [31:0] din_11_ab0;
wire [31:0] din_11_ab1;
wire [31:0] din_11_ab2;
wire [31:0] din_11_ab3;
wire [31:0] din_11_ab0_1sc;
wire [31:0] din_11_ab1_1sc;
wire [31:0] din_11_ab2_1sc;
wire [31:0] din_11_ab3_1sc;
wire [23:0] din_11_msk_ab0;
wire [23:0] din_11_msk_ab1;
wire [23:0] din_11_msk_ab2;
wire [23:0] din_11_msk_ab3;
wire [23:0] din_11_msk_ab0_1sc;
wire [23:0] din_11_msk_ab1_1sc;
wire [23:0] din_11_msk_ab2_1sc;
wire [23:0] din_11_msk_ab3_1sc;
wire [31:0] din_12_ab0;
wire [31:0] din_12_ab1;
wire [31:0] din_12_ab2;
wire [31:0] din_12_ab3;
wire [31:0] din_12_ab0_1sc;
wire [31:0] din_12_ab1_1sc;
wire [31:0] din_12_ab2_1sc;
wire [31:0] din_12_ab3_1sc;
wire [23:0] din_12_msk_ab0;
wire [23:0] din_12_msk_ab1;
wire [23:0] din_12_msk_ab2;
wire [23:0] din_12_msk_ab3;
wire [23:0] din_12_msk_ab0_1sc;
wire [23:0] din_12_msk_ab1_1sc;
wire [23:0] din_12_msk_ab2_1sc;
wire [23:0] din_12_msk_ab3_1sc;
wire [31:0] din_13_ab0;
wire [31:0] din_13_ab1;
wire [31:0] din_13_ab2;
wire [31:0] din_13_ab3;
wire [31:0] din_13_ab0_1sc;
wire [31:0] din_13_ab1_1sc;
wire [31:0] din_13_ab2_1sc;
wire [31:0] din_13_ab3_1sc;
wire [23:0] din_13_msk_ab0;
wire [23:0] din_13_msk_ab1;
wire [23:0] din_13_msk_ab2;
wire [23:0] din_13_msk_ab3;
wire [23:0] din_13_msk_ab0_1sc;
wire [23:0] din_13_msk_ab1_1sc;
wire [23:0] din_13_msk_ab2_1sc;
wire [23:0] din_13_msk_ab3_1sc;
wire [31:0] din_14_ab0;
wire [31:0] din_14_ab1;
wire [31:0] din_14_ab2;
wire [31:0] din_14_ab3;
wire [31:0] din_14_ab0_1sc;
wire [31:0] din_14_ab1_1sc;
wire [31:0] din_14_ab2_1sc;
wire [31:0] din_14_ab3_1sc;
wire [23:0] din_14_msk_ab0;
wire [23:0] din_14_msk_ab1;
wire [23:0] din_14_msk_ab2;
wire [23:0] din_14_msk_ab3;
wire [23:0] din_14_msk_ab0_1sc;
wire [23:0] din_14_msk_ab1_1sc;
wire [23:0] din_14_msk_ab2_1sc;
wire [23:0] din_14_msk_ab3_1sc;
wire [31:0] din_15_ab0;
wire [31:0] din_15_ab1;
wire [31:0] din_15_ab2;
wire [31:0] din_15_ab3;
wire [31:0] din_15_ab0_1sc;
wire [31:0] din_15_ab1_1sc;
wire [31:0] din_15_ab2_1sc;
wire [31:0] din_15_ab3_1sc;
wire [23:0] din_15_msk_ab0;
wire [23:0] din_15_msk_ab1;
wire [23:0] din_15_msk_ab2;
wire [23:0] din_15_msk_ab3;
wire [23:0] din_15_msk_ab0_1sc;
wire [23:0] din_15_msk_ab1_1sc;
wire [23:0] din_15_msk_ab2_1sc;
wire [23:0] din_15_msk_ab3_1sc;
wire [31:0] din_16_ab0;
wire [31:0] din_16_ab1;
wire [31:0] din_16_ab2;
wire [31:0] din_16_ab3;
wire [31:0] din_16_ab0_1sc;
wire [31:0] din_16_ab1_1sc;
wire [31:0] din_16_ab2_1sc;
wire [31:0] din_16_ab3_1sc;
wire [23:0] din_16_msk_ab0;
wire [23:0] din_16_msk_ab1;
wire [23:0] din_16_msk_ab2;
wire [23:0] din_16_msk_ab3;
wire [23:0] din_16_msk_ab0_1sc;
wire [23:0] din_16_msk_ab1_1sc;
wire [23:0] din_16_msk_ab2_1sc;
wire [23:0] din_16_msk_ab3_1sc;
wire [31:0] din_17_ab0;
wire [31:0] din_17_ab1;
wire [31:0] din_17_ab2;
wire [31:0] din_17_ab3;
wire [31:0] din_17_ab0_1sc;
wire [31:0] din_17_ab1_1sc;
wire [31:0] din_17_ab2_1sc;
wire [31:0] din_17_ab3_1sc;
wire [23:0] din_17_msk_ab0;
wire [23:0] din_17_msk_ab1;
wire [23:0] din_17_msk_ab2;
wire [23:0] din_17_msk_ab3;
wire [23:0] din_17_msk_ab0_1sc;
wire [23:0] din_17_msk_ab1_1sc;
wire [23:0] din_17_msk_ab2_1sc;
wire [23:0] din_17_msk_ab3_1sc;
wire [31:0] din_18_ab0;
wire [31:0] din_18_ab1;
wire [31:0] din_18_ab2;
wire [31:0] din_18_ab3;
wire [31:0] din_18_ab0_1sc;
wire [31:0] din_18_ab1_1sc;
wire [31:0] din_18_ab2_1sc;
wire [31:0] din_18_ab3_1sc;
wire [23:0] din_18_msk_ab0;
wire [23:0] din_18_msk_ab1;
wire [23:0] din_18_msk_ab2;
wire [23:0] din_18_msk_ab3;
wire [23:0] din_18_msk_ab0_1sc;
wire [23:0] din_18_msk_ab1_1sc;
wire [23:0] din_18_msk_ab2_1sc;
wire [23:0] din_18_msk_ab3_1sc;
wire [31:0] din_19_ab0;
wire [31:0] din_19_ab1;
wire [31:0] din_19_ab2;
wire [31:0] din_19_ab3;
wire [31:0] din_19_ab0_1sc;
wire [31:0] din_19_ab1_1sc;
wire [31:0] din_19_ab2_1sc;
wire [31:0] din_19_ab3_1sc;
wire [23:0] din_19_msk_ab0;
wire [23:0] din_19_msk_ab1;
wire [23:0] din_19_msk_ab2;
wire [23:0] din_19_msk_ab3;
wire [23:0] din_19_msk_ab0_1sc;
wire [23:0] din_19_msk_ab1_1sc;
wire [23:0] din_19_msk_ab2_1sc;
wire [23:0] din_19_msk_ab3_1sc;
wire [31:0] din_20_ab0;
wire [31:0] din_20_ab1;
wire [31:0] din_20_ab2;
wire [31:0] din_20_ab3;
wire [31:0] din_20_ab0_1sc;
wire [31:0] din_20_ab1_1sc;
wire [31:0] din_20_ab2_1sc;
wire [31:0] din_20_ab3_1sc;
wire [23:0] din_20_msk_ab0;
wire [23:0] din_20_msk_ab1;
wire [23:0] din_20_msk_ab2;
wire [23:0] din_20_msk_ab3;
wire [23:0] din_20_msk_ab0_1sc;
wire [23:0] din_20_msk_ab1_1sc;
wire [23:0] din_20_msk_ab2_1sc;
wire [23:0] din_20_msk_ab3_1sc;
wire [31:0] din_21_ab0;
wire [31:0] din_21_ab1;
wire [31:0] din_21_ab2;
wire [31:0] din_21_ab3;
wire [31:0] din_21_ab0_1sc;
wire [31:0] din_21_ab1_1sc;
wire [31:0] din_21_ab2_1sc;
wire [31:0] din_21_ab3_1sc;
wire [23:0] din_21_msk_ab0;
wire [23:0] din_21_msk_ab1;
wire [23:0] din_21_msk_ab2;
wire [23:0] din_21_msk_ab3;
wire [23:0] din_21_msk_ab0_1sc;
wire [23:0] din_21_msk_ab1_1sc;
wire [23:0] din_21_msk_ab2_1sc;
wire [23:0] din_21_msk_ab3_1sc;
wire [31:0] din_22_ab0;
wire [31:0] din_22_ab1;
wire [31:0] din_22_ab2;
wire [31:0] din_22_ab3;
wire [31:0] din_22_ab0_1sc;
wire [31:0] din_22_ab1_1sc;
wire [31:0] din_22_ab2_1sc;
wire [31:0] din_22_ab3_1sc;
wire [23:0] din_22_msk_ab0;
wire [23:0] din_22_msk_ab1;
wire [23:0] din_22_msk_ab2;
wire [23:0] din_22_msk_ab3;
wire [23:0] din_22_msk_ab0_1sc;
wire [23:0] din_22_msk_ab1_1sc;
wire [23:0] din_22_msk_ab2_1sc;
wire [23:0] din_22_msk_ab3_1sc;
wire [31:0] din_23_ab0;
wire [31:0] din_23_ab1;
wire [31:0] din_23_ab2;
wire [31:0] din_23_ab3;
wire [31:0] din_23_ab0_1sc;
wire [31:0] din_23_ab1_1sc;
wire [31:0] din_23_ab2_1sc;
wire [31:0] din_23_ab3_1sc;
wire [23:0] din_23_msk_ab0;
wire [23:0] din_23_msk_ab1;
wire [23:0] din_23_msk_ab2;
wire [23:0] din_23_msk_ab3;
wire [23:0] din_23_msk_ab0_1sc;
wire [23:0] din_23_msk_ab1_1sc;
wire [23:0] din_23_msk_ab2_1sc;
wire [23:0] din_23_msk_ab3_1sc;
wire [31:0] din_24_ab0;
wire [31:0] din_24_ab1;
wire [31:0] din_24_ab2;
wire [31:0] din_24_ab3;
wire [31:0] din_24_ab0_1sc;
wire [31:0] din_24_ab1_1sc;
wire [31:0] din_24_ab2_1sc;
wire [31:0] din_24_ab3_1sc;
wire [23:0] din_24_msk_ab0;
wire [23:0] din_24_msk_ab1;
wire [23:0] din_24_msk_ab2;
wire [23:0] din_24_msk_ab3;
wire [23:0] din_24_msk_ab0_1sc;
wire [23:0] din_24_msk_ab1_1sc;
wire [23:0] din_24_msk_ab2_1sc;
wire [23:0] din_24_msk_ab3_1sc;
wire [31:0] din_25_ab0;
wire [31:0] din_25_ab1;
wire [31:0] din_25_ab2;
wire [31:0] din_25_ab3;
wire [31:0] din_25_ab0_1sc;
wire [31:0] din_25_ab1_1sc;
wire [31:0] din_25_ab2_1sc;
wire [31:0] din_25_ab3_1sc;
wire [23:0] din_25_msk_ab0;
wire [23:0] din_25_msk_ab1;
wire [23:0] din_25_msk_ab2;
wire [23:0] din_25_msk_ab3;
wire [23:0] din_25_msk_ab0_1sc;
wire [23:0] din_25_msk_ab1_1sc;
wire [23:0] din_25_msk_ab2_1sc;
wire [23:0] din_25_msk_ab3_1sc;
wire [31:0] din_26_ab0;
wire [31:0] din_26_ab1;
wire [31:0] din_26_ab2;
wire [31:0] din_26_ab3;
wire [31:0] din_26_ab0_1sc;
wire [31:0] din_26_ab1_1sc;
wire [31:0] din_26_ab2_1sc;
wire [31:0] din_26_ab3_1sc;
wire [23:0] din_26_msk_ab0;
wire [23:0] din_26_msk_ab1;
wire [23:0] din_26_msk_ab2;
wire [23:0] din_26_msk_ab3;
wire [23:0] din_26_msk_ab0_1sc;
wire [23:0] din_26_msk_ab1_1sc;
wire [23:0] din_26_msk_ab2_1sc;
wire [23:0] din_26_msk_ab3_1sc;
wire [31:0] din_27_ab0;
wire [31:0] din_27_ab1;
wire [31:0] din_27_ab2;
wire [31:0] din_27_ab3;
wire [31:0] din_27_ab0_1sc;
wire [31:0] din_27_ab1_1sc;
wire [31:0] din_27_ab2_1sc;
wire [31:0] din_27_ab3_1sc;
wire [23:0] din_27_msk_ab0;
wire [23:0] din_27_msk_ab1;
wire [23:0] din_27_msk_ab2;
wire [23:0] din_27_msk_ab3;
wire [23:0] din_27_msk_ab0_1sc;
wire [23:0] din_27_msk_ab1_1sc;
wire [23:0] din_27_msk_ab2_1sc;
wire [23:0] din_27_msk_ab3_1sc;
wire [31:0] din_28_ab0;
wire [31:0] din_28_ab1;
wire [31:0] din_28_ab2;
wire [31:0] din_28_ab3;
wire [31:0] din_28_ab0_1sc;
wire [31:0] din_28_ab1_1sc;
wire [31:0] din_28_ab2_1sc;
wire [31:0] din_28_ab3_1sc;
wire [23:0] din_28_msk_ab0;
wire [23:0] din_28_msk_ab1;
wire [23:0] din_28_msk_ab2;
wire [23:0] din_28_msk_ab3;
wire [23:0] din_28_msk_ab0_1sc;
wire [23:0] din_28_msk_ab1_1sc;
wire [23:0] din_28_msk_ab2_1sc;
wire [23:0] din_28_msk_ab3_1sc;
wire [31:0] din_29_ab0;
wire [31:0] din_29_ab1;
wire [31:0] din_29_ab2;
wire [31:0] din_29_ab3;
wire [31:0] din_29_ab0_1sc;
wire [31:0] din_29_ab1_1sc;
wire [31:0] din_29_ab2_1sc;
wire [31:0] din_29_ab3_1sc;
wire [23:0] din_29_msk_ab0;
wire [23:0] din_29_msk_ab1;
wire [23:0] din_29_msk_ab2;
wire [23:0] din_29_msk_ab3;
wire [23:0] din_29_msk_ab0_1sc;
wire [23:0] din_29_msk_ab1_1sc;
wire [23:0] din_29_msk_ab2_1sc;
wire [23:0] din_29_msk_ab3_1sc;
wire [31:0] din_30_ab0;
wire [31:0] din_30_ab1;
wire [31:0] din_30_ab2;
wire [31:0] din_30_ab3;
wire [31:0] din_30_ab0_1sc;
wire [31:0] din_30_ab1_1sc;
wire [31:0] din_30_ab2_1sc;
wire [31:0] din_30_ab3_1sc;
wire [23:0] din_30_msk_ab0;
wire [23:0] din_30_msk_ab1;
wire [23:0] din_30_msk_ab2;
wire [23:0] din_30_msk_ab3;
wire [23:0] din_30_msk_ab0_1sc;
wire [23:0] din_30_msk_ab1_1sc;
wire [23:0] din_30_msk_ab2_1sc;
wire [23:0] din_30_msk_ab3_1sc;
wire [31:0] din_31_ab0;
wire [31:0] din_31_ab1;
wire [31:0] din_31_ab2;
wire [31:0] din_31_ab3;
wire [31:0] din_31_ab0_1sc;
wire [31:0] din_31_ab1_1sc;
wire [31:0] din_31_ab2_1sc;
wire [31:0] din_31_ab3_1sc;
wire [23:0] din_31_msk_ab0;
wire [23:0] din_31_msk_ab1;
wire [23:0] din_31_msk_ab2;
wire [23:0] din_31_msk_ab3;
wire [23:0] din_31_msk_ab0_1sc;
wire [23:0] din_31_msk_ab1_1sc;
wire [23:0] din_31_msk_ab2_1sc;
wire [23:0] din_31_msk_ab3_1sc;
wire [31:0] din_32_ab0;
wire [31:0] din_32_ab1;
wire [31:0] din_32_ab2;
wire [31:0] din_32_ab3;
wire [31:0] din_32_ab0_1sc;
wire [31:0] din_32_ab1_1sc;
wire [31:0] din_32_ab2_1sc;
wire [31:0] din_32_ab3_1sc;
wire [23:0] din_32_msk_ab0;
wire [23:0] din_32_msk_ab1;
wire [23:0] din_32_msk_ab2;
wire [23:0] din_32_msk_ab3;
wire [23:0] din_32_msk_ab0_1sc;
wire [23:0] din_32_msk_ab1_1sc;
wire [23:0] din_32_msk_ab2_1sc;
wire [23:0] din_32_msk_ab3_1sc;
wire [31:0] din_33_ab0;
wire [31:0] din_33_ab1;
wire [31:0] din_33_ab2;
wire [31:0] din_33_ab3;
wire [31:0] din_33_ab0_1sc;
wire [31:0] din_33_ab1_1sc;
wire [31:0] din_33_ab2_1sc;
wire [31:0] din_33_ab3_1sc;
wire [23:0] din_33_msk_ab0;
wire [23:0] din_33_msk_ab1;
wire [23:0] din_33_msk_ab2;
wire [23:0] din_33_msk_ab3;
wire [23:0] din_33_msk_ab0_1sc;
wire [23:0] din_33_msk_ab1_1sc;
wire [23:0] din_33_msk_ab2_1sc;
wire [23:0] din_33_msk_ab3_1sc;
wire [31:0] din_34_ab0;
wire [31:0] din_34_ab1;
wire [31:0] din_34_ab2;
wire [31:0] din_34_ab3;
wire [31:0] din_34_ab0_1sc;
wire [31:0] din_34_ab1_1sc;
wire [31:0] din_34_ab2_1sc;
wire [31:0] din_34_ab3_1sc;
wire [23:0] din_34_msk_ab0;
wire [23:0] din_34_msk_ab1;
wire [23:0] din_34_msk_ab2;
wire [23:0] din_34_msk_ab3;
wire [23:0] din_34_msk_ab0_1sc;
wire [23:0] din_34_msk_ab1_1sc;
wire [23:0] din_34_msk_ab2_1sc;
wire [23:0] din_34_msk_ab3_1sc;
wire [31:0] din_35_ab0;
wire [31:0] din_35_ab1;
wire [31:0] din_35_ab2;
wire [31:0] din_35_ab3;
wire [31:0] din_35_ab0_1sc;
wire [31:0] din_35_ab1_1sc;
wire [31:0] din_35_ab2_1sc;
wire [31:0] din_35_ab3_1sc;
wire [23:0] din_35_msk_ab0;
wire [23:0] din_35_msk_ab1;
wire [23:0] din_35_msk_ab2;
wire [23:0] din_35_msk_ab3;
wire [23:0] din_35_msk_ab0_1sc;
wire [23:0] din_35_msk_ab1_1sc;
wire [23:0] din_35_msk_ab2_1sc;
wire [23:0] din_35_msk_ab3_1sc;
wire [31:0] din_36_ab0;
wire [31:0] din_36_ab1;
wire [31:0] din_36_ab2;
wire [31:0] din_36_ab3;
wire [31:0] din_36_ab0_1sc;
wire [31:0] din_36_ab1_1sc;
wire [31:0] din_36_ab2_1sc;
wire [31:0] din_36_ab3_1sc;
wire [23:0] din_36_msk_ab0;
wire [23:0] din_36_msk_ab1;
wire [23:0] din_36_msk_ab2;
wire [23:0] din_36_msk_ab3;
wire [23:0] din_36_msk_ab0_1sc;
wire [23:0] din_36_msk_ab1_1sc;
wire [23:0] din_36_msk_ab2_1sc;
wire [23:0] din_36_msk_ab3_1sc;
wire [31:0] din_37_ab0;
wire [31:0] din_37_ab1;
wire [31:0] din_37_ab2;
wire [31:0] din_37_ab3;
wire [31:0] din_37_ab0_1sc;
wire [31:0] din_37_ab1_1sc;
wire [31:0] din_37_ab2_1sc;
wire [31:0] din_37_ab3_1sc;
wire [23:0] din_37_msk_ab0;
wire [23:0] din_37_msk_ab1;
wire [23:0] din_37_msk_ab2;
wire [23:0] din_37_msk_ab3;
wire [23:0] din_37_msk_ab0_1sc;
wire [23:0] din_37_msk_ab1_1sc;
wire [23:0] din_37_msk_ab2_1sc;
wire [23:0] din_37_msk_ab3_1sc;
wire [31:0] din_38_ab0;
wire [31:0] din_38_ab1;
wire [31:0] din_38_ab2;
wire [31:0] din_38_ab3;
wire [31:0] din_38_ab0_1sc;
wire [31:0] din_38_ab1_1sc;
wire [31:0] din_38_ab2_1sc;
wire [31:0] din_38_ab3_1sc;
wire [23:0] din_38_msk_ab0;
wire [23:0] din_38_msk_ab1;
wire [23:0] din_38_msk_ab2;
wire [23:0] din_38_msk_ab3;
wire [23:0] din_38_msk_ab0_1sc;
wire [23:0] din_38_msk_ab1_1sc;
wire [23:0] din_38_msk_ab2_1sc;
wire [23:0] din_38_msk_ab3_1sc;

assign din_signs[0] = din[0*8+7];
assign din_signs[1] = din[1*8+7];
assign din_signs[2] = din[2*8+7];
assign din_signs[3] = din[3*8+7];
assign din_signs[4] = din[4*8+7];
assign din_signs[5] = din[5*8+7];
assign din_signs[6] = din[6*8+7];
assign din_signs[7] = din[7*8+7];
assign din_signs[8] = din[8*8+7];
assign din_signs[9] = din[9*8+7];
assign din_signs[10] = din[10*8+7];
assign din_signs[11] = din[11*8+7];
assign din_signs[12] = din[12*8+7];
assign din_signs[13] = din[13*8+7];
assign din_signs[14] = din[14*8+7];
assign din_signs[15] = din[15*8+7];
assign din_signs[16] = din[16*8+7];
assign din_signs[17] = din[17*8+7];
assign din_signs[18] = din[18*8+7];
assign din_signs[19] = din[19*8+7];
assign din_signs[20] = din[20*8+7];
assign din_signs[21] = din[21*8+7];
assign din_signs[22] = din[22*8+7];
assign din_signs[23] = din[23*8+7];
assign din_signs[24] = din[24*8+7];
assign din_signs[25] = din[25*8+7];
assign din_signs[26] = din[26*8+7];
assign din_signs[27] = din[27*8+7];
assign din_signs[28] = din[28*8+7];
assign din_signs[29] = din[29*8+7];
assign din_signs[30] = din[30*8+7];
assign din_signs[31] = din[31*8+7];

hyper_pipe #(.NUM_PIPES(6),.WIDTH(32)) sign_bits_pipe (
    .clk(clk),.din(din_signs),.dout(din_signs_reg));

assign padded_din = {din[32*8-1:0], din_reg[63:8]};

mul_hash din_0_mul_hash (
    .clk(clk),
    .a(padded_din[0*8+:16]), 
    .ab0(din_0_ab0),                 
    .ab1(din_0_ab1), 
    .ab2(din_0_ab2),                 
    .ab3(din_0_ab3),
    .ab0_1sc(din_0_ab0_1sc),         
    .ab1_1sc(din_0_ab1_1sc), 
    .ab2_1sc(din_0_ab2_1sc),         
    .ab3_1sc(din_0_ab3_1sc),
    .msk_ab0(din_0_msk_ab0),        
    .msk_ab1(din_0_msk_ab1), 
    .msk_ab2(din_0_msk_ab2),        
    .msk_ab3(din_0_msk_ab3),
    .msk_ab0_1sc(din_0_msk_ab0_1sc), 
    .msk_ab1_1sc(din_0_msk_ab1_1sc), 
    .msk_ab2_1sc(din_0_msk_ab2_1sc), 
    .msk_ab3_1sc(din_0_msk_ab3_1sc)
);

mul_hash din_1_mul_hash (
    .clk(clk),
    .a(padded_din[1*8+:16]), 
    .ab0(din_1_ab0),                 
    .ab1(din_1_ab1), 
    .ab2(din_1_ab2),                 
    .ab3(din_1_ab3),
    .ab0_1sc(din_1_ab0_1sc),         
    .ab1_1sc(din_1_ab1_1sc), 
    .ab2_1sc(din_1_ab2_1sc),         
    .ab3_1sc(din_1_ab3_1sc),
    .msk_ab0(din_1_msk_ab0),        
    .msk_ab1(din_1_msk_ab1), 
    .msk_ab2(din_1_msk_ab2),        
    .msk_ab3(din_1_msk_ab3),
    .msk_ab0_1sc(din_1_msk_ab0_1sc), 
    .msk_ab1_1sc(din_1_msk_ab1_1sc), 
    .msk_ab2_1sc(din_1_msk_ab2_1sc), 
    .msk_ab3_1sc(din_1_msk_ab3_1sc)
);

mul_hash din_2_mul_hash (
    .clk(clk),
    .a(padded_din[2*8+:16]), 
    .ab0(din_2_ab0),                 
    .ab1(din_2_ab1), 
    .ab2(din_2_ab2),                 
    .ab3(din_2_ab3),
    .ab0_1sc(din_2_ab0_1sc),         
    .ab1_1sc(din_2_ab1_1sc), 
    .ab2_1sc(din_2_ab2_1sc),         
    .ab3_1sc(din_2_ab3_1sc),
    .msk_ab0(din_2_msk_ab0),        
    .msk_ab1(din_2_msk_ab1), 
    .msk_ab2(din_2_msk_ab2),        
    .msk_ab3(din_2_msk_ab3),
    .msk_ab0_1sc(din_2_msk_ab0_1sc), 
    .msk_ab1_1sc(din_2_msk_ab1_1sc), 
    .msk_ab2_1sc(din_2_msk_ab2_1sc), 
    .msk_ab3_1sc(din_2_msk_ab3_1sc)
);

mul_hash din_3_mul_hash (
    .clk(clk),
    .a(padded_din[3*8+:16]), 
    .ab0(din_3_ab0),                 
    .ab1(din_3_ab1), 
    .ab2(din_3_ab2),                 
    .ab3(din_3_ab3),
    .ab0_1sc(din_3_ab0_1sc),         
    .ab1_1sc(din_3_ab1_1sc), 
    .ab2_1sc(din_3_ab2_1sc),         
    .ab3_1sc(din_3_ab3_1sc),
    .msk_ab0(din_3_msk_ab0),        
    .msk_ab1(din_3_msk_ab1), 
    .msk_ab2(din_3_msk_ab2),        
    .msk_ab3(din_3_msk_ab3),
    .msk_ab0_1sc(din_3_msk_ab0_1sc), 
    .msk_ab1_1sc(din_3_msk_ab1_1sc), 
    .msk_ab2_1sc(din_3_msk_ab2_1sc), 
    .msk_ab3_1sc(din_3_msk_ab3_1sc)
);

mul_hash din_4_mul_hash (
    .clk(clk),
    .a(padded_din[4*8+:16]), 
    .ab0(din_4_ab0),                 
    .ab1(din_4_ab1), 
    .ab2(din_4_ab2),                 
    .ab3(din_4_ab3),
    .ab0_1sc(din_4_ab0_1sc),         
    .ab1_1sc(din_4_ab1_1sc), 
    .ab2_1sc(din_4_ab2_1sc),         
    .ab3_1sc(din_4_ab3_1sc),
    .msk_ab0(din_4_msk_ab0),        
    .msk_ab1(din_4_msk_ab1), 
    .msk_ab2(din_4_msk_ab2),        
    .msk_ab3(din_4_msk_ab3),
    .msk_ab0_1sc(din_4_msk_ab0_1sc), 
    .msk_ab1_1sc(din_4_msk_ab1_1sc), 
    .msk_ab2_1sc(din_4_msk_ab2_1sc), 
    .msk_ab3_1sc(din_4_msk_ab3_1sc)
);

mul_hash din_5_mul_hash (
    .clk(clk),
    .a(padded_din[5*8+:16]), 
    .ab0(din_5_ab0),                 
    .ab1(din_5_ab1), 
    .ab2(din_5_ab2),                 
    .ab3(din_5_ab3),
    .ab0_1sc(din_5_ab0_1sc),         
    .ab1_1sc(din_5_ab1_1sc), 
    .ab2_1sc(din_5_ab2_1sc),         
    .ab3_1sc(din_5_ab3_1sc),
    .msk_ab0(din_5_msk_ab0),        
    .msk_ab1(din_5_msk_ab1), 
    .msk_ab2(din_5_msk_ab2),        
    .msk_ab3(din_5_msk_ab3),
    .msk_ab0_1sc(din_5_msk_ab0_1sc), 
    .msk_ab1_1sc(din_5_msk_ab1_1sc), 
    .msk_ab2_1sc(din_5_msk_ab2_1sc), 
    .msk_ab3_1sc(din_5_msk_ab3_1sc)
);

mul_hash din_6_mul_hash (
    .clk(clk),
    .a(padded_din[6*8+:16]), 
    .ab0(din_6_ab0),                 
    .ab1(din_6_ab1), 
    .ab2(din_6_ab2),                 
    .ab3(din_6_ab3),
    .ab0_1sc(din_6_ab0_1sc),         
    .ab1_1sc(din_6_ab1_1sc), 
    .ab2_1sc(din_6_ab2_1sc),         
    .ab3_1sc(din_6_ab3_1sc),
    .msk_ab0(din_6_msk_ab0),        
    .msk_ab1(din_6_msk_ab1), 
    .msk_ab2(din_6_msk_ab2),        
    .msk_ab3(din_6_msk_ab3),
    .msk_ab0_1sc(din_6_msk_ab0_1sc), 
    .msk_ab1_1sc(din_6_msk_ab1_1sc), 
    .msk_ab2_1sc(din_6_msk_ab2_1sc), 
    .msk_ab3_1sc(din_6_msk_ab3_1sc)
);

mul_hash din_7_mul_hash (
    .clk(clk),
    .a(padded_din[7*8+:16]), 
    .ab0(din_7_ab0),                 
    .ab1(din_7_ab1), 
    .ab2(din_7_ab2),                 
    .ab3(din_7_ab3),
    .ab0_1sc(din_7_ab0_1sc),         
    .ab1_1sc(din_7_ab1_1sc), 
    .ab2_1sc(din_7_ab2_1sc),         
    .ab3_1sc(din_7_ab3_1sc),
    .msk_ab0(din_7_msk_ab0),        
    .msk_ab1(din_7_msk_ab1), 
    .msk_ab2(din_7_msk_ab2),        
    .msk_ab3(din_7_msk_ab3),
    .msk_ab0_1sc(din_7_msk_ab0_1sc), 
    .msk_ab1_1sc(din_7_msk_ab1_1sc), 
    .msk_ab2_1sc(din_7_msk_ab2_1sc), 
    .msk_ab3_1sc(din_7_msk_ab3_1sc)
);

mul_hash din_8_mul_hash (
    .clk(clk),
    .a(padded_din[8*8+:16]), 
    .ab0(din_8_ab0),                 
    .ab1(din_8_ab1), 
    .ab2(din_8_ab2),                 
    .ab3(din_8_ab3),
    .ab0_1sc(din_8_ab0_1sc),         
    .ab1_1sc(din_8_ab1_1sc), 
    .ab2_1sc(din_8_ab2_1sc),         
    .ab3_1sc(din_8_ab3_1sc),
    .msk_ab0(din_8_msk_ab0),        
    .msk_ab1(din_8_msk_ab1), 
    .msk_ab2(din_8_msk_ab2),        
    .msk_ab3(din_8_msk_ab3),
    .msk_ab0_1sc(din_8_msk_ab0_1sc), 
    .msk_ab1_1sc(din_8_msk_ab1_1sc), 
    .msk_ab2_1sc(din_8_msk_ab2_1sc), 
    .msk_ab3_1sc(din_8_msk_ab3_1sc)
);

mul_hash din_9_mul_hash (
    .clk(clk),
    .a(padded_din[9*8+:16]), 
    .ab0(din_9_ab0),                 
    .ab1(din_9_ab1), 
    .ab2(din_9_ab2),                 
    .ab3(din_9_ab3),
    .ab0_1sc(din_9_ab0_1sc),         
    .ab1_1sc(din_9_ab1_1sc), 
    .ab2_1sc(din_9_ab2_1sc),         
    .ab3_1sc(din_9_ab3_1sc),
    .msk_ab0(din_9_msk_ab0),        
    .msk_ab1(din_9_msk_ab1), 
    .msk_ab2(din_9_msk_ab2),        
    .msk_ab3(din_9_msk_ab3),
    .msk_ab0_1sc(din_9_msk_ab0_1sc), 
    .msk_ab1_1sc(din_9_msk_ab1_1sc), 
    .msk_ab2_1sc(din_9_msk_ab2_1sc), 
    .msk_ab3_1sc(din_9_msk_ab3_1sc)
);

mul_hash din_10_mul_hash (
    .clk(clk),
    .a(padded_din[10*8+:16]), 
    .ab0(din_10_ab0),                 
    .ab1(din_10_ab1), 
    .ab2(din_10_ab2),                 
    .ab3(din_10_ab3),
    .ab0_1sc(din_10_ab0_1sc),         
    .ab1_1sc(din_10_ab1_1sc), 
    .ab2_1sc(din_10_ab2_1sc),         
    .ab3_1sc(din_10_ab3_1sc),
    .msk_ab0(din_10_msk_ab0),        
    .msk_ab1(din_10_msk_ab1), 
    .msk_ab2(din_10_msk_ab2),        
    .msk_ab3(din_10_msk_ab3),
    .msk_ab0_1sc(din_10_msk_ab0_1sc), 
    .msk_ab1_1sc(din_10_msk_ab1_1sc), 
    .msk_ab2_1sc(din_10_msk_ab2_1sc), 
    .msk_ab3_1sc(din_10_msk_ab3_1sc)
);

mul_hash din_11_mul_hash (
    .clk(clk),
    .a(padded_din[11*8+:16]), 
    .ab0(din_11_ab0),                 
    .ab1(din_11_ab1), 
    .ab2(din_11_ab2),                 
    .ab3(din_11_ab3),
    .ab0_1sc(din_11_ab0_1sc),         
    .ab1_1sc(din_11_ab1_1sc), 
    .ab2_1sc(din_11_ab2_1sc),         
    .ab3_1sc(din_11_ab3_1sc),
    .msk_ab0(din_11_msk_ab0),        
    .msk_ab1(din_11_msk_ab1), 
    .msk_ab2(din_11_msk_ab2),        
    .msk_ab3(din_11_msk_ab3),
    .msk_ab0_1sc(din_11_msk_ab0_1sc), 
    .msk_ab1_1sc(din_11_msk_ab1_1sc), 
    .msk_ab2_1sc(din_11_msk_ab2_1sc), 
    .msk_ab3_1sc(din_11_msk_ab3_1sc)
);

mul_hash din_12_mul_hash (
    .clk(clk),
    .a(padded_din[12*8+:16]), 
    .ab0(din_12_ab0),                 
    .ab1(din_12_ab1), 
    .ab2(din_12_ab2),                 
    .ab3(din_12_ab3),
    .ab0_1sc(din_12_ab0_1sc),         
    .ab1_1sc(din_12_ab1_1sc), 
    .ab2_1sc(din_12_ab2_1sc),         
    .ab3_1sc(din_12_ab3_1sc),
    .msk_ab0(din_12_msk_ab0),        
    .msk_ab1(din_12_msk_ab1), 
    .msk_ab2(din_12_msk_ab2),        
    .msk_ab3(din_12_msk_ab3),
    .msk_ab0_1sc(din_12_msk_ab0_1sc), 
    .msk_ab1_1sc(din_12_msk_ab1_1sc), 
    .msk_ab2_1sc(din_12_msk_ab2_1sc), 
    .msk_ab3_1sc(din_12_msk_ab3_1sc)
);

mul_hash din_13_mul_hash (
    .clk(clk),
    .a(padded_din[13*8+:16]), 
    .ab0(din_13_ab0),                 
    .ab1(din_13_ab1), 
    .ab2(din_13_ab2),                 
    .ab3(din_13_ab3),
    .ab0_1sc(din_13_ab0_1sc),         
    .ab1_1sc(din_13_ab1_1sc), 
    .ab2_1sc(din_13_ab2_1sc),         
    .ab3_1sc(din_13_ab3_1sc),
    .msk_ab0(din_13_msk_ab0),        
    .msk_ab1(din_13_msk_ab1), 
    .msk_ab2(din_13_msk_ab2),        
    .msk_ab3(din_13_msk_ab3),
    .msk_ab0_1sc(din_13_msk_ab0_1sc), 
    .msk_ab1_1sc(din_13_msk_ab1_1sc), 
    .msk_ab2_1sc(din_13_msk_ab2_1sc), 
    .msk_ab3_1sc(din_13_msk_ab3_1sc)
);

mul_hash din_14_mul_hash (
    .clk(clk),
    .a(padded_din[14*8+:16]), 
    .ab0(din_14_ab0),                 
    .ab1(din_14_ab1), 
    .ab2(din_14_ab2),                 
    .ab3(din_14_ab3),
    .ab0_1sc(din_14_ab0_1sc),         
    .ab1_1sc(din_14_ab1_1sc), 
    .ab2_1sc(din_14_ab2_1sc),         
    .ab3_1sc(din_14_ab3_1sc),
    .msk_ab0(din_14_msk_ab0),        
    .msk_ab1(din_14_msk_ab1), 
    .msk_ab2(din_14_msk_ab2),        
    .msk_ab3(din_14_msk_ab3),
    .msk_ab0_1sc(din_14_msk_ab0_1sc), 
    .msk_ab1_1sc(din_14_msk_ab1_1sc), 
    .msk_ab2_1sc(din_14_msk_ab2_1sc), 
    .msk_ab3_1sc(din_14_msk_ab3_1sc)
);

mul_hash din_15_mul_hash (
    .clk(clk),
    .a(padded_din[15*8+:16]), 
    .ab0(din_15_ab0),                 
    .ab1(din_15_ab1), 
    .ab2(din_15_ab2),                 
    .ab3(din_15_ab3),
    .ab0_1sc(din_15_ab0_1sc),         
    .ab1_1sc(din_15_ab1_1sc), 
    .ab2_1sc(din_15_ab2_1sc),         
    .ab3_1sc(din_15_ab3_1sc),
    .msk_ab0(din_15_msk_ab0),        
    .msk_ab1(din_15_msk_ab1), 
    .msk_ab2(din_15_msk_ab2),        
    .msk_ab3(din_15_msk_ab3),
    .msk_ab0_1sc(din_15_msk_ab0_1sc), 
    .msk_ab1_1sc(din_15_msk_ab1_1sc), 
    .msk_ab2_1sc(din_15_msk_ab2_1sc), 
    .msk_ab3_1sc(din_15_msk_ab3_1sc)
);

mul_hash din_16_mul_hash (
    .clk(clk),
    .a(padded_din[16*8+:16]), 
    .ab0(din_16_ab0),                 
    .ab1(din_16_ab1), 
    .ab2(din_16_ab2),                 
    .ab3(din_16_ab3),
    .ab0_1sc(din_16_ab0_1sc),         
    .ab1_1sc(din_16_ab1_1sc), 
    .ab2_1sc(din_16_ab2_1sc),         
    .ab3_1sc(din_16_ab3_1sc),
    .msk_ab0(din_16_msk_ab0),        
    .msk_ab1(din_16_msk_ab1), 
    .msk_ab2(din_16_msk_ab2),        
    .msk_ab3(din_16_msk_ab3),
    .msk_ab0_1sc(din_16_msk_ab0_1sc), 
    .msk_ab1_1sc(din_16_msk_ab1_1sc), 
    .msk_ab2_1sc(din_16_msk_ab2_1sc), 
    .msk_ab3_1sc(din_16_msk_ab3_1sc)
);

mul_hash din_17_mul_hash (
    .clk(clk),
    .a(padded_din[17*8+:16]), 
    .ab0(din_17_ab0),                 
    .ab1(din_17_ab1), 
    .ab2(din_17_ab2),                 
    .ab3(din_17_ab3),
    .ab0_1sc(din_17_ab0_1sc),         
    .ab1_1sc(din_17_ab1_1sc), 
    .ab2_1sc(din_17_ab2_1sc),         
    .ab3_1sc(din_17_ab3_1sc),
    .msk_ab0(din_17_msk_ab0),        
    .msk_ab1(din_17_msk_ab1), 
    .msk_ab2(din_17_msk_ab2),        
    .msk_ab3(din_17_msk_ab3),
    .msk_ab0_1sc(din_17_msk_ab0_1sc), 
    .msk_ab1_1sc(din_17_msk_ab1_1sc), 
    .msk_ab2_1sc(din_17_msk_ab2_1sc), 
    .msk_ab3_1sc(din_17_msk_ab3_1sc)
);

mul_hash din_18_mul_hash (
    .clk(clk),
    .a(padded_din[18*8+:16]), 
    .ab0(din_18_ab0),                 
    .ab1(din_18_ab1), 
    .ab2(din_18_ab2),                 
    .ab3(din_18_ab3),
    .ab0_1sc(din_18_ab0_1sc),         
    .ab1_1sc(din_18_ab1_1sc), 
    .ab2_1sc(din_18_ab2_1sc),         
    .ab3_1sc(din_18_ab3_1sc),
    .msk_ab0(din_18_msk_ab0),        
    .msk_ab1(din_18_msk_ab1), 
    .msk_ab2(din_18_msk_ab2),        
    .msk_ab3(din_18_msk_ab3),
    .msk_ab0_1sc(din_18_msk_ab0_1sc), 
    .msk_ab1_1sc(din_18_msk_ab1_1sc), 
    .msk_ab2_1sc(din_18_msk_ab2_1sc), 
    .msk_ab3_1sc(din_18_msk_ab3_1sc)
);

mul_hash din_19_mul_hash (
    .clk(clk),
    .a(padded_din[19*8+:16]), 
    .ab0(din_19_ab0),                 
    .ab1(din_19_ab1), 
    .ab2(din_19_ab2),                 
    .ab3(din_19_ab3),
    .ab0_1sc(din_19_ab0_1sc),         
    .ab1_1sc(din_19_ab1_1sc), 
    .ab2_1sc(din_19_ab2_1sc),         
    .ab3_1sc(din_19_ab3_1sc),
    .msk_ab0(din_19_msk_ab0),        
    .msk_ab1(din_19_msk_ab1), 
    .msk_ab2(din_19_msk_ab2),        
    .msk_ab3(din_19_msk_ab3),
    .msk_ab0_1sc(din_19_msk_ab0_1sc), 
    .msk_ab1_1sc(din_19_msk_ab1_1sc), 
    .msk_ab2_1sc(din_19_msk_ab2_1sc), 
    .msk_ab3_1sc(din_19_msk_ab3_1sc)
);

mul_hash din_20_mul_hash (
    .clk(clk),
    .a(padded_din[20*8+:16]), 
    .ab0(din_20_ab0),                 
    .ab1(din_20_ab1), 
    .ab2(din_20_ab2),                 
    .ab3(din_20_ab3),
    .ab0_1sc(din_20_ab0_1sc),         
    .ab1_1sc(din_20_ab1_1sc), 
    .ab2_1sc(din_20_ab2_1sc),         
    .ab3_1sc(din_20_ab3_1sc),
    .msk_ab0(din_20_msk_ab0),        
    .msk_ab1(din_20_msk_ab1), 
    .msk_ab2(din_20_msk_ab2),        
    .msk_ab3(din_20_msk_ab3),
    .msk_ab0_1sc(din_20_msk_ab0_1sc), 
    .msk_ab1_1sc(din_20_msk_ab1_1sc), 
    .msk_ab2_1sc(din_20_msk_ab2_1sc), 
    .msk_ab3_1sc(din_20_msk_ab3_1sc)
);

mul_hash din_21_mul_hash (
    .clk(clk),
    .a(padded_din[21*8+:16]), 
    .ab0(din_21_ab0),                 
    .ab1(din_21_ab1), 
    .ab2(din_21_ab2),                 
    .ab3(din_21_ab3),
    .ab0_1sc(din_21_ab0_1sc),         
    .ab1_1sc(din_21_ab1_1sc), 
    .ab2_1sc(din_21_ab2_1sc),         
    .ab3_1sc(din_21_ab3_1sc),
    .msk_ab0(din_21_msk_ab0),        
    .msk_ab1(din_21_msk_ab1), 
    .msk_ab2(din_21_msk_ab2),        
    .msk_ab3(din_21_msk_ab3),
    .msk_ab0_1sc(din_21_msk_ab0_1sc), 
    .msk_ab1_1sc(din_21_msk_ab1_1sc), 
    .msk_ab2_1sc(din_21_msk_ab2_1sc), 
    .msk_ab3_1sc(din_21_msk_ab3_1sc)
);

mul_hash din_22_mul_hash (
    .clk(clk),
    .a(padded_din[22*8+:16]), 
    .ab0(din_22_ab0),                 
    .ab1(din_22_ab1), 
    .ab2(din_22_ab2),                 
    .ab3(din_22_ab3),
    .ab0_1sc(din_22_ab0_1sc),         
    .ab1_1sc(din_22_ab1_1sc), 
    .ab2_1sc(din_22_ab2_1sc),         
    .ab3_1sc(din_22_ab3_1sc),
    .msk_ab0(din_22_msk_ab0),        
    .msk_ab1(din_22_msk_ab1), 
    .msk_ab2(din_22_msk_ab2),        
    .msk_ab3(din_22_msk_ab3),
    .msk_ab0_1sc(din_22_msk_ab0_1sc), 
    .msk_ab1_1sc(din_22_msk_ab1_1sc), 
    .msk_ab2_1sc(din_22_msk_ab2_1sc), 
    .msk_ab3_1sc(din_22_msk_ab3_1sc)
);

mul_hash din_23_mul_hash (
    .clk(clk),
    .a(padded_din[23*8+:16]), 
    .ab0(din_23_ab0),                 
    .ab1(din_23_ab1), 
    .ab2(din_23_ab2),                 
    .ab3(din_23_ab3),
    .ab0_1sc(din_23_ab0_1sc),         
    .ab1_1sc(din_23_ab1_1sc), 
    .ab2_1sc(din_23_ab2_1sc),         
    .ab3_1sc(din_23_ab3_1sc),
    .msk_ab0(din_23_msk_ab0),        
    .msk_ab1(din_23_msk_ab1), 
    .msk_ab2(din_23_msk_ab2),        
    .msk_ab3(din_23_msk_ab3),
    .msk_ab0_1sc(din_23_msk_ab0_1sc), 
    .msk_ab1_1sc(din_23_msk_ab1_1sc), 
    .msk_ab2_1sc(din_23_msk_ab2_1sc), 
    .msk_ab3_1sc(din_23_msk_ab3_1sc)
);

mul_hash din_24_mul_hash (
    .clk(clk),
    .a(padded_din[24*8+:16]), 
    .ab0(din_24_ab0),                 
    .ab1(din_24_ab1), 
    .ab2(din_24_ab2),                 
    .ab3(din_24_ab3),
    .ab0_1sc(din_24_ab0_1sc),         
    .ab1_1sc(din_24_ab1_1sc), 
    .ab2_1sc(din_24_ab2_1sc),         
    .ab3_1sc(din_24_ab3_1sc),
    .msk_ab0(din_24_msk_ab0),        
    .msk_ab1(din_24_msk_ab1), 
    .msk_ab2(din_24_msk_ab2),        
    .msk_ab3(din_24_msk_ab3),
    .msk_ab0_1sc(din_24_msk_ab0_1sc), 
    .msk_ab1_1sc(din_24_msk_ab1_1sc), 
    .msk_ab2_1sc(din_24_msk_ab2_1sc), 
    .msk_ab3_1sc(din_24_msk_ab3_1sc)
);

mul_hash din_25_mul_hash (
    .clk(clk),
    .a(padded_din[25*8+:16]), 
    .ab0(din_25_ab0),                 
    .ab1(din_25_ab1), 
    .ab2(din_25_ab2),                 
    .ab3(din_25_ab3),
    .ab0_1sc(din_25_ab0_1sc),         
    .ab1_1sc(din_25_ab1_1sc), 
    .ab2_1sc(din_25_ab2_1sc),         
    .ab3_1sc(din_25_ab3_1sc),
    .msk_ab0(din_25_msk_ab0),        
    .msk_ab1(din_25_msk_ab1), 
    .msk_ab2(din_25_msk_ab2),        
    .msk_ab3(din_25_msk_ab3),
    .msk_ab0_1sc(din_25_msk_ab0_1sc), 
    .msk_ab1_1sc(din_25_msk_ab1_1sc), 
    .msk_ab2_1sc(din_25_msk_ab2_1sc), 
    .msk_ab3_1sc(din_25_msk_ab3_1sc)
);

mul_hash din_26_mul_hash (
    .clk(clk),
    .a(padded_din[26*8+:16]), 
    .ab0(din_26_ab0),                 
    .ab1(din_26_ab1), 
    .ab2(din_26_ab2),                 
    .ab3(din_26_ab3),
    .ab0_1sc(din_26_ab0_1sc),         
    .ab1_1sc(din_26_ab1_1sc), 
    .ab2_1sc(din_26_ab2_1sc),         
    .ab3_1sc(din_26_ab3_1sc),
    .msk_ab0(din_26_msk_ab0),        
    .msk_ab1(din_26_msk_ab1), 
    .msk_ab2(din_26_msk_ab2),        
    .msk_ab3(din_26_msk_ab3),
    .msk_ab0_1sc(din_26_msk_ab0_1sc), 
    .msk_ab1_1sc(din_26_msk_ab1_1sc), 
    .msk_ab2_1sc(din_26_msk_ab2_1sc), 
    .msk_ab3_1sc(din_26_msk_ab3_1sc)
);

mul_hash din_27_mul_hash (
    .clk(clk),
    .a(padded_din[27*8+:16]), 
    .ab0(din_27_ab0),                 
    .ab1(din_27_ab1), 
    .ab2(din_27_ab2),                 
    .ab3(din_27_ab3),
    .ab0_1sc(din_27_ab0_1sc),         
    .ab1_1sc(din_27_ab1_1sc), 
    .ab2_1sc(din_27_ab2_1sc),         
    .ab3_1sc(din_27_ab3_1sc),
    .msk_ab0(din_27_msk_ab0),        
    .msk_ab1(din_27_msk_ab1), 
    .msk_ab2(din_27_msk_ab2),        
    .msk_ab3(din_27_msk_ab3),
    .msk_ab0_1sc(din_27_msk_ab0_1sc), 
    .msk_ab1_1sc(din_27_msk_ab1_1sc), 
    .msk_ab2_1sc(din_27_msk_ab2_1sc), 
    .msk_ab3_1sc(din_27_msk_ab3_1sc)
);

mul_hash din_28_mul_hash (
    .clk(clk),
    .a(padded_din[28*8+:16]), 
    .ab0(din_28_ab0),                 
    .ab1(din_28_ab1), 
    .ab2(din_28_ab2),                 
    .ab3(din_28_ab3),
    .ab0_1sc(din_28_ab0_1sc),         
    .ab1_1sc(din_28_ab1_1sc), 
    .ab2_1sc(din_28_ab2_1sc),         
    .ab3_1sc(din_28_ab3_1sc),
    .msk_ab0(din_28_msk_ab0),        
    .msk_ab1(din_28_msk_ab1), 
    .msk_ab2(din_28_msk_ab2),        
    .msk_ab3(din_28_msk_ab3),
    .msk_ab0_1sc(din_28_msk_ab0_1sc), 
    .msk_ab1_1sc(din_28_msk_ab1_1sc), 
    .msk_ab2_1sc(din_28_msk_ab2_1sc), 
    .msk_ab3_1sc(din_28_msk_ab3_1sc)
);

mul_hash din_29_mul_hash (
    .clk(clk),
    .a(padded_din[29*8+:16]), 
    .ab0(din_29_ab0),                 
    .ab1(din_29_ab1), 
    .ab2(din_29_ab2),                 
    .ab3(din_29_ab3),
    .ab0_1sc(din_29_ab0_1sc),         
    .ab1_1sc(din_29_ab1_1sc), 
    .ab2_1sc(din_29_ab2_1sc),         
    .ab3_1sc(din_29_ab3_1sc),
    .msk_ab0(din_29_msk_ab0),        
    .msk_ab1(din_29_msk_ab1), 
    .msk_ab2(din_29_msk_ab2),        
    .msk_ab3(din_29_msk_ab3),
    .msk_ab0_1sc(din_29_msk_ab0_1sc), 
    .msk_ab1_1sc(din_29_msk_ab1_1sc), 
    .msk_ab2_1sc(din_29_msk_ab2_1sc), 
    .msk_ab3_1sc(din_29_msk_ab3_1sc)
);

mul_hash din_30_mul_hash (
    .clk(clk),
    .a(padded_din[30*8+:16]), 
    .ab0(din_30_ab0),                 
    .ab1(din_30_ab1), 
    .ab2(din_30_ab2),                 
    .ab3(din_30_ab3),
    .ab0_1sc(din_30_ab0_1sc),         
    .ab1_1sc(din_30_ab1_1sc), 
    .ab2_1sc(din_30_ab2_1sc),         
    .ab3_1sc(din_30_ab3_1sc),
    .msk_ab0(din_30_msk_ab0),        
    .msk_ab1(din_30_msk_ab1), 
    .msk_ab2(din_30_msk_ab2),        
    .msk_ab3(din_30_msk_ab3),
    .msk_ab0_1sc(din_30_msk_ab0_1sc), 
    .msk_ab1_1sc(din_30_msk_ab1_1sc), 
    .msk_ab2_1sc(din_30_msk_ab2_1sc), 
    .msk_ab3_1sc(din_30_msk_ab3_1sc)
);

mul_hash din_31_mul_hash (
    .clk(clk),
    .a(padded_din[31*8+:16]), 
    .ab0(din_31_ab0),                 
    .ab1(din_31_ab1), 
    .ab2(din_31_ab2),                 
    .ab3(din_31_ab3),
    .ab0_1sc(din_31_ab0_1sc),         
    .ab1_1sc(din_31_ab1_1sc), 
    .ab2_1sc(din_31_ab2_1sc),         
    .ab3_1sc(din_31_ab3_1sc),
    .msk_ab0(din_31_msk_ab0),        
    .msk_ab1(din_31_msk_ab1), 
    .msk_ab2(din_31_msk_ab2),        
    .msk_ab3(din_31_msk_ab3),
    .msk_ab0_1sc(din_31_msk_ab0_1sc), 
    .msk_ab1_1sc(din_31_msk_ab1_1sc), 
    .msk_ab2_1sc(din_31_msk_ab2_1sc), 
    .msk_ab3_1sc(din_31_msk_ab3_1sc)
);

mul_hash din_32_mul_hash (
    .clk(clk),
    .a(padded_din[32*8+:16]), 
    .ab0(din_32_ab0),                 
    .ab1(din_32_ab1), 
    .ab2(din_32_ab2),                 
    .ab3(din_32_ab3),
    .ab0_1sc(din_32_ab0_1sc),         
    .ab1_1sc(din_32_ab1_1sc), 
    .ab2_1sc(din_32_ab2_1sc),         
    .ab3_1sc(din_32_ab3_1sc),
    .msk_ab0(din_32_msk_ab0),        
    .msk_ab1(din_32_msk_ab1), 
    .msk_ab2(din_32_msk_ab2),        
    .msk_ab3(din_32_msk_ab3),
    .msk_ab0_1sc(din_32_msk_ab0_1sc), 
    .msk_ab1_1sc(din_32_msk_ab1_1sc), 
    .msk_ab2_1sc(din_32_msk_ab2_1sc), 
    .msk_ab3_1sc(din_32_msk_ab3_1sc)
);

mul_hash din_33_mul_hash (
    .clk(clk),
    .a(padded_din[33*8+:16]), 
    .ab0(din_33_ab0),                 
    .ab1(din_33_ab1), 
    .ab2(din_33_ab2),                 
    .ab3(din_33_ab3),
    .ab0_1sc(din_33_ab0_1sc),         
    .ab1_1sc(din_33_ab1_1sc), 
    .ab2_1sc(din_33_ab2_1sc),         
    .ab3_1sc(din_33_ab3_1sc),
    .msk_ab0(din_33_msk_ab0),        
    .msk_ab1(din_33_msk_ab1), 
    .msk_ab2(din_33_msk_ab2),        
    .msk_ab3(din_33_msk_ab3),
    .msk_ab0_1sc(din_33_msk_ab0_1sc), 
    .msk_ab1_1sc(din_33_msk_ab1_1sc), 
    .msk_ab2_1sc(din_33_msk_ab2_1sc), 
    .msk_ab3_1sc(din_33_msk_ab3_1sc)
);

mul_hash din_34_mul_hash (
    .clk(clk),
    .a(padded_din[34*8+:16]), 
    .ab0(din_34_ab0),                 
    .ab1(din_34_ab1), 
    .ab2(din_34_ab2),                 
    .ab3(din_34_ab3),
    .ab0_1sc(din_34_ab0_1sc),         
    .ab1_1sc(din_34_ab1_1sc), 
    .ab2_1sc(din_34_ab2_1sc),         
    .ab3_1sc(din_34_ab3_1sc),
    .msk_ab0(din_34_msk_ab0),        
    .msk_ab1(din_34_msk_ab1), 
    .msk_ab2(din_34_msk_ab2),        
    .msk_ab3(din_34_msk_ab3),
    .msk_ab0_1sc(din_34_msk_ab0_1sc), 
    .msk_ab1_1sc(din_34_msk_ab1_1sc), 
    .msk_ab2_1sc(din_34_msk_ab2_1sc), 
    .msk_ab3_1sc(din_34_msk_ab3_1sc)
);

mul_hash din_35_mul_hash (
    .clk(clk),
    .a(padded_din[35*8+:16]), 
    .ab0(din_35_ab0),                 
    .ab1(din_35_ab1), 
    .ab2(din_35_ab2),                 
    .ab3(din_35_ab3),
    .ab0_1sc(din_35_ab0_1sc),         
    .ab1_1sc(din_35_ab1_1sc), 
    .ab2_1sc(din_35_ab2_1sc),         
    .ab3_1sc(din_35_ab3_1sc),
    .msk_ab0(din_35_msk_ab0),        
    .msk_ab1(din_35_msk_ab1), 
    .msk_ab2(din_35_msk_ab2),        
    .msk_ab3(din_35_msk_ab3),
    .msk_ab0_1sc(din_35_msk_ab0_1sc), 
    .msk_ab1_1sc(din_35_msk_ab1_1sc), 
    .msk_ab2_1sc(din_35_msk_ab2_1sc), 
    .msk_ab3_1sc(din_35_msk_ab3_1sc)
);

mul_hash din_36_mul_hash (
    .clk(clk),
    .a(padded_din[36*8+:16]), 
    .ab0(din_36_ab0),                 
    .ab1(din_36_ab1), 
    .ab2(din_36_ab2),                 
    .ab3(din_36_ab3),
    .ab0_1sc(din_36_ab0_1sc),         
    .ab1_1sc(din_36_ab1_1sc), 
    .ab2_1sc(din_36_ab2_1sc),         
    .ab3_1sc(din_36_ab3_1sc),
    .msk_ab0(din_36_msk_ab0),        
    .msk_ab1(din_36_msk_ab1), 
    .msk_ab2(din_36_msk_ab2),        
    .msk_ab3(din_36_msk_ab3),
    .msk_ab0_1sc(din_36_msk_ab0_1sc), 
    .msk_ab1_1sc(din_36_msk_ab1_1sc), 
    .msk_ab2_1sc(din_36_msk_ab2_1sc), 
    .msk_ab3_1sc(din_36_msk_ab3_1sc)
);

mul_hash din_37_mul_hash (
    .clk(clk),
    .a(padded_din[37*8+:16]), 
    .ab0(din_37_ab0),                 
    .ab1(din_37_ab1), 
    .ab2(din_37_ab2),                 
    .ab3(din_37_ab3),
    .ab0_1sc(din_37_ab0_1sc),         
    .ab1_1sc(din_37_ab1_1sc), 
    .ab2_1sc(din_37_ab2_1sc),         
    .ab3_1sc(din_37_ab3_1sc),
    .msk_ab0(din_37_msk_ab0),        
    .msk_ab1(din_37_msk_ab1), 
    .msk_ab2(din_37_msk_ab2),        
    .msk_ab3(din_37_msk_ab3),
    .msk_ab0_1sc(din_37_msk_ab0_1sc), 
    .msk_ab1_1sc(din_37_msk_ab1_1sc), 
    .msk_ab2_1sc(din_37_msk_ab2_1sc), 
    .msk_ab3_1sc(din_37_msk_ab3_1sc)
);

mul_hash din_38_mul_hash (
    .clk(clk),
    .a(padded_din[38*8+:16]), 
    .ab0(din_38_ab0),                 
    .ab1(din_38_ab1), 
    .ab2(din_38_ab2),                 
    .ab3(din_38_ab3),
    .ab0_1sc(din_38_ab0_1sc),         
    .ab1_1sc(din_38_ab1_1sc), 
    .ab2_1sc(din_38_ab2_1sc),         
    .ab3_1sc(din_38_ab3_1sc),
    .msk_ab0(din_38_msk_ab0),        
    .msk_ab1(din_38_msk_ab1), 
    .msk_ab2(din_38_msk_ab2),        
    .msk_ab3(din_38_msk_ab3),
    .msk_ab0_1sc(din_38_msk_ab0_1sc), 
    .msk_ab1_1sc(din_38_msk_ab1_1sc), 
    .msk_ab2_1sc(din_38_msk_ab2_1sc), 
    .msk_ab3_1sc(din_38_msk_ab3_1sc)
);


//Valid signals
assign din_valid_0_0 = din_valid & din_valid_reg;
assign din_valid_1_0 = din_valid & din_valid_reg;
assign din_valid_0_1 = din_valid & din_valid_reg;
assign din_valid_1_1 = din_valid & din_valid_reg;
assign din_valid_0_2 = din_valid & din_valid_reg;
assign din_valid_1_2 = din_valid & din_valid_reg;
assign din_valid_0_3 = din_valid & din_valid_reg;
assign din_valid_1_3 = din_valid & din_valid_reg;
assign din_valid_0_4 = din_valid & din_valid_reg;
assign din_valid_1_4 = din_valid & din_valid_reg;
assign din_valid_0_5 = din_valid & din_valid_reg;
assign din_valid_1_5 = din_valid & din_valid_reg;
assign din_valid_0_6 = din_valid & din_valid_reg;
assign din_valid_1_6 = din_valid & din_valid_reg;
assign din_valid_0_7 = din_valid;
assign din_valid_1_7 = din_valid;
assign din_valid_0_8 = din_valid;
assign din_valid_1_8 = din_valid;
assign din_valid_0_9 = din_valid;
assign din_valid_1_9 = din_valid;
assign din_valid_0_10 = din_valid;
assign din_valid_1_10 = din_valid;
assign din_valid_0_11 = din_valid;
assign din_valid_1_11 = din_valid;
assign din_valid_0_12 = din_valid;
assign din_valid_1_12 = din_valid;
assign din_valid_0_13 = din_valid;
assign din_valid_1_13 = din_valid;
assign din_valid_0_14 = din_valid;
assign din_valid_1_14 = din_valid;
assign din_valid_0_15 = din_valid;
assign din_valid_1_15 = din_valid;
assign din_valid_0_16 = din_valid;
assign din_valid_1_16 = din_valid;
assign din_valid_0_17 = din_valid;
assign din_valid_1_17 = din_valid;
assign din_valid_0_18 = din_valid;
assign din_valid_1_18 = din_valid;
assign din_valid_0_19 = din_valid;
assign din_valid_1_19 = din_valid;
assign din_valid_0_20 = din_valid;
assign din_valid_1_20 = din_valid;
assign din_valid_0_21 = din_valid;
assign din_valid_1_21 = din_valid;
assign din_valid_0_22 = din_valid;
assign din_valid_1_22 = din_valid;
assign din_valid_0_23 = din_valid;
assign din_valid_1_23 = din_valid;
assign din_valid_0_24 = din_valid;
assign din_valid_1_24 = din_valid;
assign din_valid_0_25 = din_valid;
assign din_valid_1_25 = din_valid;
assign din_valid_0_26 = din_valid;
assign din_valid_1_26 = din_valid;
assign din_valid_0_27 = din_valid;
assign din_valid_1_27 = din_valid;
assign din_valid_0_28 = din_valid;
assign din_valid_1_28 = din_valid;
assign din_valid_0_29 = din_valid;
assign din_valid_1_29 = din_valid;
assign din_valid_0_30 = din_valid;
assign din_valid_1_30 = din_valid;
assign din_valid_0_31 = din_valid;
assign din_valid_1_31 = din_valid;

assign din_valid_2_0 = din_valid & din_valid_reg;
assign din_valid_2_1 = din_valid & din_valid_reg;
assign din_valid_2_2 = din_valid & din_valid_reg;
assign din_valid_2_3 = din_valid & din_valid_reg;
assign din_valid_2_4 = din_valid & din_valid_reg;
assign din_valid_2_5 = din_valid & din_valid_reg;
assign din_valid_2_6 = din_valid;
assign din_valid_2_7 = din_valid;
assign din_valid_2_8 = din_valid;
assign din_valid_2_9 = din_valid;
assign din_valid_2_10 = din_valid;
assign din_valid_2_11 = din_valid;
assign din_valid_2_12 = din_valid;
assign din_valid_2_13 = din_valid;
assign din_valid_2_14 = din_valid;
assign din_valid_2_15 = din_valid;
assign din_valid_2_16 = din_valid;
assign din_valid_2_17 = din_valid;
assign din_valid_2_18 = din_valid;
assign din_valid_2_19 = din_valid;
assign din_valid_2_20 = din_valid;
assign din_valid_2_21 = din_valid;
assign din_valid_2_22 = din_valid;
assign din_valid_2_23 = din_valid;
assign din_valid_2_24 = din_valid;
assign din_valid_2_25 = din_valid;
assign din_valid_2_26 = din_valid;
assign din_valid_2_27 = din_valid;
assign din_valid_2_28 = din_valid;
assign din_valid_2_29 = din_valid;
assign din_valid_2_30 = din_valid;
assign din_valid_2_31 = din_valid;

assign din_valid_3_0 = din_valid & din_valid_reg;
assign din_valid_3_1 = din_valid & din_valid_reg;
assign din_valid_3_2 = din_valid & din_valid_reg;
assign din_valid_3_3 = din_valid & din_valid_reg;
assign din_valid_3_4 = din_valid & din_valid_reg;
assign din_valid_3_5 = din_valid;
assign din_valid_3_6 = din_valid;
assign din_valid_3_7 = din_valid;
assign din_valid_3_8 = din_valid;
assign din_valid_3_9 = din_valid;
assign din_valid_3_10 = din_valid;
assign din_valid_3_11 = din_valid;
assign din_valid_3_12 = din_valid;
assign din_valid_3_13 = din_valid;
assign din_valid_3_14 = din_valid;
assign din_valid_3_15 = din_valid;
assign din_valid_3_16 = din_valid;
assign din_valid_3_17 = din_valid;
assign din_valid_3_18 = din_valid;
assign din_valid_3_19 = din_valid;
assign din_valid_3_20 = din_valid;
assign din_valid_3_21 = din_valid;
assign din_valid_3_22 = din_valid;
assign din_valid_3_23 = din_valid;
assign din_valid_3_24 = din_valid;
assign din_valid_3_25 = din_valid;
assign din_valid_3_26 = din_valid;
assign din_valid_3_27 = din_valid;
assign din_valid_3_28 = din_valid;
assign din_valid_3_29 = din_valid;
assign din_valid_3_30 = din_valid;
assign din_valid_3_31 = din_valid;

assign din_valid_4_0 = din_valid & din_valid_reg;
assign din_valid_4_1 = din_valid & din_valid_reg;
assign din_valid_4_2 = din_valid & din_valid_reg;
assign din_valid_4_3 = din_valid & din_valid_reg;
assign din_valid_4_4 = din_valid;
assign din_valid_4_5 = din_valid;
assign din_valid_4_6 = din_valid;
assign din_valid_4_7 = din_valid;
assign din_valid_4_8 = din_valid;
assign din_valid_4_9 = din_valid;
assign din_valid_4_10 = din_valid;
assign din_valid_4_11 = din_valid;
assign din_valid_4_12 = din_valid;
assign din_valid_4_13 = din_valid;
assign din_valid_4_14 = din_valid;
assign din_valid_4_15 = din_valid;
assign din_valid_4_16 = din_valid;
assign din_valid_4_17 = din_valid;
assign din_valid_4_18 = din_valid;
assign din_valid_4_19 = din_valid;
assign din_valid_4_20 = din_valid;
assign din_valid_4_21 = din_valid;
assign din_valid_4_22 = din_valid;
assign din_valid_4_23 = din_valid;
assign din_valid_4_24 = din_valid;
assign din_valid_4_25 = din_valid;
assign din_valid_4_26 = din_valid;
assign din_valid_4_27 = din_valid;
assign din_valid_4_28 = din_valid;
assign din_valid_4_29 = din_valid;
assign din_valid_4_30 = din_valid;
assign din_valid_4_31 = din_valid;

assign din_valid_5_0 = din_valid & din_valid_reg;
assign din_valid_5_1 = din_valid & din_valid_reg;
assign din_valid_5_2 = din_valid & din_valid_reg;
assign din_valid_5_3 = din_valid;
assign din_valid_5_4 = din_valid;
assign din_valid_5_5 = din_valid;
assign din_valid_5_6 = din_valid;
assign din_valid_5_7 = din_valid;
assign din_valid_5_8 = din_valid;
assign din_valid_5_9 = din_valid;
assign din_valid_5_10 = din_valid;
assign din_valid_5_11 = din_valid;
assign din_valid_5_12 = din_valid;
assign din_valid_5_13 = din_valid;
assign din_valid_5_14 = din_valid;
assign din_valid_5_15 = din_valid;
assign din_valid_5_16 = din_valid;
assign din_valid_5_17 = din_valid;
assign din_valid_5_18 = din_valid;
assign din_valid_5_19 = din_valid;
assign din_valid_5_20 = din_valid;
assign din_valid_5_21 = din_valid;
assign din_valid_5_22 = din_valid;
assign din_valid_5_23 = din_valid;
assign din_valid_5_24 = din_valid;
assign din_valid_5_25 = din_valid;
assign din_valid_5_26 = din_valid;
assign din_valid_5_27 = din_valid;
assign din_valid_5_28 = din_valid;
assign din_valid_5_29 = din_valid;
assign din_valid_5_30 = din_valid;
assign din_valid_5_31 = din_valid;

assign din_valid_6_0 = din_valid & din_valid_reg;
assign din_valid_6_1 = din_valid & din_valid_reg;
assign din_valid_6_2 = din_valid;
assign din_valid_6_3 = din_valid;
assign din_valid_6_4 = din_valid;
assign din_valid_6_5 = din_valid;
assign din_valid_6_6 = din_valid;
assign din_valid_6_7 = din_valid;
assign din_valid_6_8 = din_valid;
assign din_valid_6_9 = din_valid;
assign din_valid_6_10 = din_valid;
assign din_valid_6_11 = din_valid;
assign din_valid_6_12 = din_valid;
assign din_valid_6_13 = din_valid;
assign din_valid_6_14 = din_valid;
assign din_valid_6_15 = din_valid;
assign din_valid_6_16 = din_valid;
assign din_valid_6_17 = din_valid;
assign din_valid_6_18 = din_valid;
assign din_valid_6_19 = din_valid;
assign din_valid_6_20 = din_valid;
assign din_valid_6_21 = din_valid;
assign din_valid_6_22 = din_valid;
assign din_valid_6_23 = din_valid;
assign din_valid_6_24 = din_valid;
assign din_valid_6_25 = din_valid;
assign din_valid_6_26 = din_valid;
assign din_valid_6_27 = din_valid;
assign din_valid_6_28 = din_valid;
assign din_valid_6_29 = din_valid;
assign din_valid_6_30 = din_valid;
assign din_valid_6_31 = din_valid;

assign din_valid_7_0 = din_valid & din_valid_reg;
assign din_valid_7_1 = din_valid;
assign din_valid_7_2 = din_valid;
assign din_valid_7_3 = din_valid;
assign din_valid_7_4 = din_valid;
assign din_valid_7_5 = din_valid;
assign din_valid_7_6 = din_valid;
assign din_valid_7_7 = din_valid;
assign din_valid_7_8 = din_valid;
assign din_valid_7_9 = din_valid;
assign din_valid_7_10 = din_valid;
assign din_valid_7_11 = din_valid;
assign din_valid_7_12 = din_valid;
assign din_valid_7_13 = din_valid;
assign din_valid_7_14 = din_valid;
assign din_valid_7_15 = din_valid;
assign din_valid_7_16 = din_valid;
assign din_valid_7_17 = din_valid;
assign din_valid_7_18 = din_valid;
assign din_valid_7_19 = din_valid;
assign din_valid_7_20 = din_valid;
assign din_valid_7_21 = din_valid;
assign din_valid_7_22 = din_valid;
assign din_valid_7_23 = din_valid;
assign din_valid_7_24 = din_valid;
assign din_valid_7_25 = din_valid;
assign din_valid_7_26 = din_valid;
assign din_valid_7_27 = din_valid;
assign din_valid_7_28 = din_valid;
assign din_valid_7_29 = din_valid;
assign din_valid_7_30 = din_valid;
assign din_valid_7_31 = din_valid;


always @ (posedge clk) begin
    //din_reg <= din[127:64];
    din_reg <= din[255:192];
    // din_reg <= din[63:0];
    din_valid_reg <= din_valid;
end

hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_0_pipe (
    .clk(clk),.din(din_valid_0_0),.dout(addr_valid_0_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_1_pipe (
    .clk(clk),.din(din_valid_0_1),.dout(addr_valid_0_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_2_pipe (
    .clk(clk),.din(din_valid_0_2),.dout(addr_valid_0_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_3_pipe (
    .clk(clk),.din(din_valid_0_3),.dout(addr_valid_0_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_4_pipe (
    .clk(clk),.din(din_valid_0_4),.dout(addr_valid_0_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_5_pipe (
    .clk(clk),.din(din_valid_0_5),.dout(addr_valid_0_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_6_pipe (
    .clk(clk),.din(din_valid_0_6),.dout(addr_valid_0_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_7_pipe (
    .clk(clk),.din(din_valid_0_7),.dout(addr_valid_0_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_8_pipe (
    .clk(clk),.din(din_valid_0_8),.dout(addr_valid_0_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_9_pipe (
    .clk(clk),.din(din_valid_0_9),.dout(addr_valid_0_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_10_pipe (
    .clk(clk),.din(din_valid_0_10),.dout(addr_valid_0_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_11_pipe (
    .clk(clk),.din(din_valid_0_11),.dout(addr_valid_0_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_12_pipe (
    .clk(clk),.din(din_valid_0_12),.dout(addr_valid_0_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_13_pipe (
    .clk(clk),.din(din_valid_0_13),.dout(addr_valid_0_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_14_pipe (
    .clk(clk),.din(din_valid_0_14),.dout(addr_valid_0_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_15_pipe (
    .clk(clk),.din(din_valid_0_15),.dout(addr_valid_0_15));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_16_pipe (
    .clk(clk),.din(din_valid_0_16),.dout(addr_valid_0_16));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_17_pipe (
    .clk(clk),.din(din_valid_0_17),.dout(addr_valid_0_17));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_18_pipe (
    .clk(clk),.din(din_valid_0_18),.dout(addr_valid_0_18));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_19_pipe (
    .clk(clk),.din(din_valid_0_19),.dout(addr_valid_0_19));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_20_pipe (
    .clk(clk),.din(din_valid_0_20),.dout(addr_valid_0_20));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_21_pipe (
    .clk(clk),.din(din_valid_0_21),.dout(addr_valid_0_21));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_22_pipe (
    .clk(clk),.din(din_valid_0_22),.dout(addr_valid_0_22));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_23_pipe (
    .clk(clk),.din(din_valid_0_23),.dout(addr_valid_0_23));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_24_pipe (
    .clk(clk),.din(din_valid_0_24),.dout(addr_valid_0_24));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_25_pipe (
    .clk(clk),.din(din_valid_0_25),.dout(addr_valid_0_25));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_26_pipe (
    .clk(clk),.din(din_valid_0_26),.dout(addr_valid_0_26));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_27_pipe (
    .clk(clk),.din(din_valid_0_27),.dout(addr_valid_0_27));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_28_pipe (
    .clk(clk),.din(din_valid_0_28),.dout(addr_valid_0_28));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_29_pipe (
    .clk(clk),.din(din_valid_0_29),.dout(addr_valid_0_29));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_30_pipe (
    .clk(clk),.din(din_valid_0_30),.dout(addr_valid_0_30));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_31_pipe (
    .clk(clk),.din(din_valid_0_31),.dout(addr_valid_0_31));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_0_pipe (
    .clk(clk),.din(din_valid_1_0),.dout(addr_valid_1_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_1_pipe (
    .clk(clk),.din(din_valid_1_1),.dout(addr_valid_1_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_2_pipe (
    .clk(clk),.din(din_valid_1_2),.dout(addr_valid_1_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_3_pipe (
    .clk(clk),.din(din_valid_1_3),.dout(addr_valid_1_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_4_pipe (
    .clk(clk),.din(din_valid_1_4),.dout(addr_valid_1_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_5_pipe (
    .clk(clk),.din(din_valid_1_5),.dout(addr_valid_1_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_6_pipe (
    .clk(clk),.din(din_valid_1_6),.dout(addr_valid_1_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_7_pipe (
    .clk(clk),.din(din_valid_1_7),.dout(addr_valid_1_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_8_pipe (
    .clk(clk),.din(din_valid_1_8),.dout(addr_valid_1_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_9_pipe (
    .clk(clk),.din(din_valid_1_9),.dout(addr_valid_1_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_10_pipe (
    .clk(clk),.din(din_valid_1_10),.dout(addr_valid_1_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_11_pipe (
    .clk(clk),.din(din_valid_1_11),.dout(addr_valid_1_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_12_pipe (
    .clk(clk),.din(din_valid_1_12),.dout(addr_valid_1_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_13_pipe (
    .clk(clk),.din(din_valid_1_13),.dout(addr_valid_1_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_14_pipe (
    .clk(clk),.din(din_valid_1_14),.dout(addr_valid_1_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_15_pipe (
    .clk(clk),.din(din_valid_1_15),.dout(addr_valid_1_15));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_16_pipe (
    .clk(clk),.din(din_valid_1_16),.dout(addr_valid_1_16));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_17_pipe (
    .clk(clk),.din(din_valid_1_17),.dout(addr_valid_1_17));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_18_pipe (
    .clk(clk),.din(din_valid_1_18),.dout(addr_valid_1_18));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_19_pipe (
    .clk(clk),.din(din_valid_1_19),.dout(addr_valid_1_19));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_20_pipe (
    .clk(clk),.din(din_valid_1_20),.dout(addr_valid_1_20));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_21_pipe (
    .clk(clk),.din(din_valid_1_21),.dout(addr_valid_1_21));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_22_pipe (
    .clk(clk),.din(din_valid_1_22),.dout(addr_valid_1_22));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_23_pipe (
    .clk(clk),.din(din_valid_1_23),.dout(addr_valid_1_23));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_24_pipe (
    .clk(clk),.din(din_valid_1_24),.dout(addr_valid_1_24));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_25_pipe (
    .clk(clk),.din(din_valid_1_25),.dout(addr_valid_1_25));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_26_pipe (
    .clk(clk),.din(din_valid_1_26),.dout(addr_valid_1_26));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_27_pipe (
    .clk(clk),.din(din_valid_1_27),.dout(addr_valid_1_27));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_28_pipe (
    .clk(clk),.din(din_valid_1_28),.dout(addr_valid_1_28));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_29_pipe (
    .clk(clk),.din(din_valid_1_29),.dout(addr_valid_1_29));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_30_pipe (
    .clk(clk),.din(din_valid_1_30),.dout(addr_valid_1_30));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_31_pipe (
    .clk(clk),.din(din_valid_1_31),.dout(addr_valid_1_31));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_0_pipe (
    .clk(clk),.din(din_valid_2_0),.dout(addr_valid_2_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_1_pipe (
    .clk(clk),.din(din_valid_2_1),.dout(addr_valid_2_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_2_pipe (
    .clk(clk),.din(din_valid_2_2),.dout(addr_valid_2_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_3_pipe (
    .clk(clk),.din(din_valid_2_3),.dout(addr_valid_2_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_4_pipe (
    .clk(clk),.din(din_valid_2_4),.dout(addr_valid_2_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_5_pipe (
    .clk(clk),.din(din_valid_2_5),.dout(addr_valid_2_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_6_pipe (
    .clk(clk),.din(din_valid_2_6),.dout(addr_valid_2_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_7_pipe (
    .clk(clk),.din(din_valid_2_7),.dout(addr_valid_2_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_8_pipe (
    .clk(clk),.din(din_valid_2_8),.dout(addr_valid_2_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_9_pipe (
    .clk(clk),.din(din_valid_2_9),.dout(addr_valid_2_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_10_pipe (
    .clk(clk),.din(din_valid_2_10),.dout(addr_valid_2_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_11_pipe (
    .clk(clk),.din(din_valid_2_11),.dout(addr_valid_2_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_12_pipe (
    .clk(clk),.din(din_valid_2_12),.dout(addr_valid_2_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_13_pipe (
    .clk(clk),.din(din_valid_2_13),.dout(addr_valid_2_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_14_pipe (
    .clk(clk),.din(din_valid_2_14),.dout(addr_valid_2_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_15_pipe (
    .clk(clk),.din(din_valid_2_15),.dout(addr_valid_2_15));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_16_pipe (
    .clk(clk),.din(din_valid_2_16),.dout(addr_valid_2_16));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_17_pipe (
    .clk(clk),.din(din_valid_2_17),.dout(addr_valid_2_17));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_18_pipe (
    .clk(clk),.din(din_valid_2_18),.dout(addr_valid_2_18));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_19_pipe (
    .clk(clk),.din(din_valid_2_19),.dout(addr_valid_2_19));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_20_pipe (
    .clk(clk),.din(din_valid_2_20),.dout(addr_valid_2_20));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_21_pipe (
    .clk(clk),.din(din_valid_2_21),.dout(addr_valid_2_21));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_22_pipe (
    .clk(clk),.din(din_valid_2_22),.dout(addr_valid_2_22));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_23_pipe (
    .clk(clk),.din(din_valid_2_23),.dout(addr_valid_2_23));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_24_pipe (
    .clk(clk),.din(din_valid_2_24),.dout(addr_valid_2_24));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_25_pipe (
    .clk(clk),.din(din_valid_2_25),.dout(addr_valid_2_25));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_26_pipe (
    .clk(clk),.din(din_valid_2_26),.dout(addr_valid_2_26));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_27_pipe (
    .clk(clk),.din(din_valid_2_27),.dout(addr_valid_2_27));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_28_pipe (
    .clk(clk),.din(din_valid_2_28),.dout(addr_valid_2_28));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_29_pipe (
    .clk(clk),.din(din_valid_2_29),.dout(addr_valid_2_29));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_30_pipe (
    .clk(clk),.din(din_valid_2_30),.dout(addr_valid_2_30));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_31_pipe (
    .clk(clk),.din(din_valid_2_31),.dout(addr_valid_2_31));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_0_pipe (
    .clk(clk),.din(din_valid_3_0),.dout(addr_valid_3_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_1_pipe (
    .clk(clk),.din(din_valid_3_1),.dout(addr_valid_3_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_2_pipe (
    .clk(clk),.din(din_valid_3_2),.dout(addr_valid_3_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_3_pipe (
    .clk(clk),.din(din_valid_3_3),.dout(addr_valid_3_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_4_pipe (
    .clk(clk),.din(din_valid_3_4),.dout(addr_valid_3_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_5_pipe (
    .clk(clk),.din(din_valid_3_5),.dout(addr_valid_3_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_6_pipe (
    .clk(clk),.din(din_valid_3_6),.dout(addr_valid_3_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_7_pipe (
    .clk(clk),.din(din_valid_3_7),.dout(addr_valid_3_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_8_pipe (
    .clk(clk),.din(din_valid_3_8),.dout(addr_valid_3_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_9_pipe (
    .clk(clk),.din(din_valid_3_9),.dout(addr_valid_3_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_10_pipe (
    .clk(clk),.din(din_valid_3_10),.dout(addr_valid_3_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_11_pipe (
    .clk(clk),.din(din_valid_3_11),.dout(addr_valid_3_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_12_pipe (
    .clk(clk),.din(din_valid_3_12),.dout(addr_valid_3_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_13_pipe (
    .clk(clk),.din(din_valid_3_13),.dout(addr_valid_3_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_14_pipe (
    .clk(clk),.din(din_valid_3_14),.dout(addr_valid_3_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_15_pipe (
    .clk(clk),.din(din_valid_3_15),.dout(addr_valid_3_15));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_16_pipe (
    .clk(clk),.din(din_valid_3_16),.dout(addr_valid_3_16));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_17_pipe (
    .clk(clk),.din(din_valid_3_17),.dout(addr_valid_3_17));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_18_pipe (
    .clk(clk),.din(din_valid_3_18),.dout(addr_valid_3_18));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_19_pipe (
    .clk(clk),.din(din_valid_3_19),.dout(addr_valid_3_19));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_20_pipe (
    .clk(clk),.din(din_valid_3_20),.dout(addr_valid_3_20));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_21_pipe (
    .clk(clk),.din(din_valid_3_21),.dout(addr_valid_3_21));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_22_pipe (
    .clk(clk),.din(din_valid_3_22),.dout(addr_valid_3_22));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_23_pipe (
    .clk(clk),.din(din_valid_3_23),.dout(addr_valid_3_23));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_24_pipe (
    .clk(clk),.din(din_valid_3_24),.dout(addr_valid_3_24));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_25_pipe (
    .clk(clk),.din(din_valid_3_25),.dout(addr_valid_3_25));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_26_pipe (
    .clk(clk),.din(din_valid_3_26),.dout(addr_valid_3_26));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_27_pipe (
    .clk(clk),.din(din_valid_3_27),.dout(addr_valid_3_27));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_28_pipe (
    .clk(clk),.din(din_valid_3_28),.dout(addr_valid_3_28));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_29_pipe (
    .clk(clk),.din(din_valid_3_29),.dout(addr_valid_3_29));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_30_pipe (
    .clk(clk),.din(din_valid_3_30),.dout(addr_valid_3_30));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_31_pipe (
    .clk(clk),.din(din_valid_3_31),.dout(addr_valid_3_31));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_0_pipe (
    .clk(clk),.din(din_valid_4_0),.dout(addr_valid_4_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_1_pipe (
    .clk(clk),.din(din_valid_4_1),.dout(addr_valid_4_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_2_pipe (
    .clk(clk),.din(din_valid_4_2),.dout(addr_valid_4_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_3_pipe (
    .clk(clk),.din(din_valid_4_3),.dout(addr_valid_4_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_4_pipe (
    .clk(clk),.din(din_valid_4_4),.dout(addr_valid_4_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_5_pipe (
    .clk(clk),.din(din_valid_4_5),.dout(addr_valid_4_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_6_pipe (
    .clk(clk),.din(din_valid_4_6),.dout(addr_valid_4_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_7_pipe (
    .clk(clk),.din(din_valid_4_7),.dout(addr_valid_4_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_8_pipe (
    .clk(clk),.din(din_valid_4_8),.dout(addr_valid_4_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_9_pipe (
    .clk(clk),.din(din_valid_4_9),.dout(addr_valid_4_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_10_pipe (
    .clk(clk),.din(din_valid_4_10),.dout(addr_valid_4_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_11_pipe (
    .clk(clk),.din(din_valid_4_11),.dout(addr_valid_4_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_12_pipe (
    .clk(clk),.din(din_valid_4_12),.dout(addr_valid_4_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_13_pipe (
    .clk(clk),.din(din_valid_4_13),.dout(addr_valid_4_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_14_pipe (
    .clk(clk),.din(din_valid_4_14),.dout(addr_valid_4_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_15_pipe (
    .clk(clk),.din(din_valid_4_15),.dout(addr_valid_4_15));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_16_pipe (
    .clk(clk),.din(din_valid_4_16),.dout(addr_valid_4_16));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_17_pipe (
    .clk(clk),.din(din_valid_4_17),.dout(addr_valid_4_17));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_18_pipe (
    .clk(clk),.din(din_valid_4_18),.dout(addr_valid_4_18));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_19_pipe (
    .clk(clk),.din(din_valid_4_19),.dout(addr_valid_4_19));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_20_pipe (
    .clk(clk),.din(din_valid_4_20),.dout(addr_valid_4_20));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_21_pipe (
    .clk(clk),.din(din_valid_4_21),.dout(addr_valid_4_21));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_22_pipe (
    .clk(clk),.din(din_valid_4_22),.dout(addr_valid_4_22));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_23_pipe (
    .clk(clk),.din(din_valid_4_23),.dout(addr_valid_4_23));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_24_pipe (
    .clk(clk),.din(din_valid_4_24),.dout(addr_valid_4_24));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_25_pipe (
    .clk(clk),.din(din_valid_4_25),.dout(addr_valid_4_25));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_26_pipe (
    .clk(clk),.din(din_valid_4_26),.dout(addr_valid_4_26));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_27_pipe (
    .clk(clk),.din(din_valid_4_27),.dout(addr_valid_4_27));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_28_pipe (
    .clk(clk),.din(din_valid_4_28),.dout(addr_valid_4_28));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_29_pipe (
    .clk(clk),.din(din_valid_4_29),.dout(addr_valid_4_29));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_30_pipe (
    .clk(clk),.din(din_valid_4_30),.dout(addr_valid_4_30));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_31_pipe (
    .clk(clk),.din(din_valid_4_31),.dout(addr_valid_4_31));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_0_pipe (
    .clk(clk),.din(din_valid_5_0),.dout(addr_valid_5_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_1_pipe (
    .clk(clk),.din(din_valid_5_1),.dout(addr_valid_5_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_2_pipe (
    .clk(clk),.din(din_valid_5_2),.dout(addr_valid_5_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_3_pipe (
    .clk(clk),.din(din_valid_5_3),.dout(addr_valid_5_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_4_pipe (
    .clk(clk),.din(din_valid_5_4),.dout(addr_valid_5_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_5_pipe (
    .clk(clk),.din(din_valid_5_5),.dout(addr_valid_5_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_6_pipe (
    .clk(clk),.din(din_valid_5_6),.dout(addr_valid_5_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_7_pipe (
    .clk(clk),.din(din_valid_5_7),.dout(addr_valid_5_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_8_pipe (
    .clk(clk),.din(din_valid_5_8),.dout(addr_valid_5_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_9_pipe (
    .clk(clk),.din(din_valid_5_9),.dout(addr_valid_5_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_10_pipe (
    .clk(clk),.din(din_valid_5_10),.dout(addr_valid_5_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_11_pipe (
    .clk(clk),.din(din_valid_5_11),.dout(addr_valid_5_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_12_pipe (
    .clk(clk),.din(din_valid_5_12),.dout(addr_valid_5_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_13_pipe (
    .clk(clk),.din(din_valid_5_13),.dout(addr_valid_5_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_14_pipe (
    .clk(clk),.din(din_valid_5_14),.dout(addr_valid_5_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_15_pipe (
    .clk(clk),.din(din_valid_5_15),.dout(addr_valid_5_15));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_16_pipe (
    .clk(clk),.din(din_valid_5_16),.dout(addr_valid_5_16));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_17_pipe (
    .clk(clk),.din(din_valid_5_17),.dout(addr_valid_5_17));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_18_pipe (
    .clk(clk),.din(din_valid_5_18),.dout(addr_valid_5_18));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_19_pipe (
    .clk(clk),.din(din_valid_5_19),.dout(addr_valid_5_19));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_20_pipe (
    .clk(clk),.din(din_valid_5_20),.dout(addr_valid_5_20));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_21_pipe (
    .clk(clk),.din(din_valid_5_21),.dout(addr_valid_5_21));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_22_pipe (
    .clk(clk),.din(din_valid_5_22),.dout(addr_valid_5_22));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_23_pipe (
    .clk(clk),.din(din_valid_5_23),.dout(addr_valid_5_23));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_24_pipe (
    .clk(clk),.din(din_valid_5_24),.dout(addr_valid_5_24));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_25_pipe (
    .clk(clk),.din(din_valid_5_25),.dout(addr_valid_5_25));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_26_pipe (
    .clk(clk),.din(din_valid_5_26),.dout(addr_valid_5_26));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_27_pipe (
    .clk(clk),.din(din_valid_5_27),.dout(addr_valid_5_27));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_28_pipe (
    .clk(clk),.din(din_valid_5_28),.dout(addr_valid_5_28));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_29_pipe (
    .clk(clk),.din(din_valid_5_29),.dout(addr_valid_5_29));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_30_pipe (
    .clk(clk),.din(din_valid_5_30),.dout(addr_valid_5_30));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_31_pipe (
    .clk(clk),.din(din_valid_5_31),.dout(addr_valid_5_31));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_0_pipe (
    .clk(clk),.din(din_valid_6_0),.dout(addr_valid_6_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_1_pipe (
    .clk(clk),.din(din_valid_6_1),.dout(addr_valid_6_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_2_pipe (
    .clk(clk),.din(din_valid_6_2),.dout(addr_valid_6_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_3_pipe (
    .clk(clk),.din(din_valid_6_3),.dout(addr_valid_6_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_4_pipe (
    .clk(clk),.din(din_valid_6_4),.dout(addr_valid_6_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_5_pipe (
    .clk(clk),.din(din_valid_6_5),.dout(addr_valid_6_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_6_pipe (
    .clk(clk),.din(din_valid_6_6),.dout(addr_valid_6_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_7_pipe (
    .clk(clk),.din(din_valid_6_7),.dout(addr_valid_6_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_8_pipe (
    .clk(clk),.din(din_valid_6_8),.dout(addr_valid_6_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_9_pipe (
    .clk(clk),.din(din_valid_6_9),.dout(addr_valid_6_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_10_pipe (
    .clk(clk),.din(din_valid_6_10),.dout(addr_valid_6_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_11_pipe (
    .clk(clk),.din(din_valid_6_11),.dout(addr_valid_6_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_12_pipe (
    .clk(clk),.din(din_valid_6_12),.dout(addr_valid_6_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_13_pipe (
    .clk(clk),.din(din_valid_6_13),.dout(addr_valid_6_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_14_pipe (
    .clk(clk),.din(din_valid_6_14),.dout(addr_valid_6_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_15_pipe (
    .clk(clk),.din(din_valid_6_15),.dout(addr_valid_6_15));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_16_pipe (
    .clk(clk),.din(din_valid_6_16),.dout(addr_valid_6_16));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_17_pipe (
    .clk(clk),.din(din_valid_6_17),.dout(addr_valid_6_17));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_18_pipe (
    .clk(clk),.din(din_valid_6_18),.dout(addr_valid_6_18));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_19_pipe (
    .clk(clk),.din(din_valid_6_19),.dout(addr_valid_6_19));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_20_pipe (
    .clk(clk),.din(din_valid_6_20),.dout(addr_valid_6_20));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_21_pipe (
    .clk(clk),.din(din_valid_6_21),.dout(addr_valid_6_21));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_22_pipe (
    .clk(clk),.din(din_valid_6_22),.dout(addr_valid_6_22));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_23_pipe (
    .clk(clk),.din(din_valid_6_23),.dout(addr_valid_6_23));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_24_pipe (
    .clk(clk),.din(din_valid_6_24),.dout(addr_valid_6_24));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_25_pipe (
    .clk(clk),.din(din_valid_6_25),.dout(addr_valid_6_25));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_26_pipe (
    .clk(clk),.din(din_valid_6_26),.dout(addr_valid_6_26));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_27_pipe (
    .clk(clk),.din(din_valid_6_27),.dout(addr_valid_6_27));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_28_pipe (
    .clk(clk),.din(din_valid_6_28),.dout(addr_valid_6_28));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_29_pipe (
    .clk(clk),.din(din_valid_6_29),.dout(addr_valid_6_29));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_30_pipe (
    .clk(clk),.din(din_valid_6_30),.dout(addr_valid_6_30));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_31_pipe (
    .clk(clk),.din(din_valid_6_31),.dout(addr_valid_6_31));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_0_pipe (
    .clk(clk),.din(din_valid_7_0),.dout(addr_valid_7_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_1_pipe (
    .clk(clk),.din(din_valid_7_1),.dout(addr_valid_7_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_2_pipe (
    .clk(clk),.din(din_valid_7_2),.dout(addr_valid_7_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_3_pipe (
    .clk(clk),.din(din_valid_7_3),.dout(addr_valid_7_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_4_pipe (
    .clk(clk),.din(din_valid_7_4),.dout(addr_valid_7_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_5_pipe (
    .clk(clk),.din(din_valid_7_5),.dout(addr_valid_7_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_6_pipe (
    .clk(clk),.din(din_valid_7_6),.dout(addr_valid_7_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_7_pipe (
    .clk(clk),.din(din_valid_7_7),.dout(addr_valid_7_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_8_pipe (
    .clk(clk),.din(din_valid_7_8),.dout(addr_valid_7_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_9_pipe (
    .clk(clk),.din(din_valid_7_9),.dout(addr_valid_7_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_10_pipe (
    .clk(clk),.din(din_valid_7_10),.dout(addr_valid_7_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_11_pipe (
    .clk(clk),.din(din_valid_7_11),.dout(addr_valid_7_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_12_pipe (
    .clk(clk),.din(din_valid_7_12),.dout(addr_valid_7_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_13_pipe (
    .clk(clk),.din(din_valid_7_13),.dout(addr_valid_7_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_14_pipe (
    .clk(clk),.din(din_valid_7_14),.dout(addr_valid_7_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_15_pipe (
    .clk(clk),.din(din_valid_7_15),.dout(addr_valid_7_15));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_16_pipe (
    .clk(clk),.din(din_valid_7_16),.dout(addr_valid_7_16));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_17_pipe (
    .clk(clk),.din(din_valid_7_17),.dout(addr_valid_7_17));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_18_pipe (
    .clk(clk),.din(din_valid_7_18),.dout(addr_valid_7_18));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_19_pipe (
    .clk(clk),.din(din_valid_7_19),.dout(addr_valid_7_19));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_20_pipe (
    .clk(clk),.din(din_valid_7_20),.dout(addr_valid_7_20));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_21_pipe (
    .clk(clk),.din(din_valid_7_21),.dout(addr_valid_7_21));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_22_pipe (
    .clk(clk),.din(din_valid_7_22),.dout(addr_valid_7_22));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_23_pipe (
    .clk(clk),.din(din_valid_7_23),.dout(addr_valid_7_23));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_24_pipe (
    .clk(clk),.din(din_valid_7_24),.dout(addr_valid_7_24));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_25_pipe (
    .clk(clk),.din(din_valid_7_25),.dout(addr_valid_7_25));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_26_pipe (
    .clk(clk),.din(din_valid_7_26),.dout(addr_valid_7_26));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_27_pipe (
    .clk(clk),.din(din_valid_7_27),.dout(addr_valid_7_27));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_28_pipe (
    .clk(clk),.din(din_valid_7_28),.dout(addr_valid_7_28));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_29_pipe (
    .clk(clk),.din(din_valid_7_29),.dout(addr_valid_7_29));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_30_pipe (
    .clk(clk),.din(din_valid_7_30),.dout(addr_valid_7_30));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_31_pipe (
    .clk(clk),.din(din_valid_7_31),.dout(addr_valid_7_31));

// Mask and Nbits is dependent on bucket number
// data selection is dependent on first byte location
acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_0_calc (
           .clk(clk), .sign(din_signs_reg[0]), 
           .p(addr_0_0),
           .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
           .a0b0_1sc(din_0_ab0_1sc), .a0b1_1sc(din_0_ab1_1sc), .a0b2_1sc(din_0_ab2_1sc), .a0b3_1sc(din_0_ab3_1sc),
           .msk_a0b0(din_0_msk_ab0), .msk_a0b1(din_0_msk_ab1), .msk_a0b2(din_0_msk_ab2), .msk_a0b3(din_0_msk_ab3),
           .msk_a0b0_1sc(din_0_msk_ab0_1sc), .msk_a0b1_1sc(din_0_msk_ab1_1sc), .msk_a0b2_1sc(din_0_msk_ab2_1sc), .msk_a0b3_1sc(din_0_msk_ab3_1sc),

           .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2),
           .a1b0_1sc(din_2_ab0_1sc), .a1b1_1sc(din_2_ab1_1sc), .a1b2_1sc(din_2_ab2_1sc),
           .msk_a1b0(din_2_msk_ab0), .msk_a1b1(din_2_msk_ab1), .msk_a1b2(din_2_msk_ab2),
           .msk_a1b0_1sc(din_2_msk_ab0_1sc), .msk_a1b1_1sc(din_2_msk_ab1_1sc), .msk_a1b2_1sc(din_2_msk_ab2_1sc),

           .a2b0(din_4_ab0), .a2b1(din_4_ab1),
           .a2b0_1sc(din_4_ab0_1sc), .a2b1_1sc(din_4_ab1_1sc),
           .msk_a2b0(din_4_msk_ab0), .msk_a2b1(din_4_msk_ab1),
           .msk_a2b0_1sc(din_4_msk_ab0_1sc), .msk_a2b1_1sc(din_4_msk_ab1_1sc),
           
           .a3b0(din_6_ab0),
           .a3b0_1sc(din_6_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_1_calc (
           .clk(clk), .sign(din_signs_reg[1]), 
           .p(addr_0_1),
           .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
           .a0b0_1sc(din_1_ab0_1sc), .a0b1_1sc(din_1_ab1_1sc), .a0b2_1sc(din_1_ab2_1sc), .a0b3_1sc(din_1_ab3_1sc),
           .msk_a0b0(din_1_msk_ab0), .msk_a0b1(din_1_msk_ab1), .msk_a0b2(din_1_msk_ab2), .msk_a0b3(din_1_msk_ab3),
           .msk_a0b0_1sc(din_1_msk_ab0_1sc), .msk_a0b1_1sc(din_1_msk_ab1_1sc), .msk_a0b2_1sc(din_1_msk_ab2_1sc), .msk_a0b3_1sc(din_1_msk_ab3_1sc),

           .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2),
           .a1b0_1sc(din_3_ab0_1sc), .a1b1_1sc(din_3_ab1_1sc), .a1b2_1sc(din_3_ab2_1sc),
           .msk_a1b0(din_3_msk_ab0), .msk_a1b1(din_3_msk_ab1), .msk_a1b2(din_3_msk_ab2),
           .msk_a1b0_1sc(din_3_msk_ab0_1sc), .msk_a1b1_1sc(din_3_msk_ab1_1sc), .msk_a1b2_1sc(din_3_msk_ab2_1sc),

           .a2b0(din_5_ab0), .a2b1(din_5_ab1),
           .a2b0_1sc(din_5_ab0_1sc), .a2b1_1sc(din_5_ab1_1sc),
           .msk_a2b0(din_5_msk_ab0), .msk_a2b1(din_5_msk_ab1),
           .msk_a2b0_1sc(din_5_msk_ab0_1sc), .msk_a2b1_1sc(din_5_msk_ab1_1sc),
           
           .a3b0(din_7_ab0),
           .a3b0_1sc(din_7_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_2_calc (
           .clk(clk), .sign(din_signs_reg[2]), 
           .p(addr_0_2),
           .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
           .a0b0_1sc(din_2_ab0_1sc), .a0b1_1sc(din_2_ab1_1sc), .a0b2_1sc(din_2_ab2_1sc), .a0b3_1sc(din_2_ab3_1sc),
           .msk_a0b0(din_2_msk_ab0), .msk_a0b1(din_2_msk_ab1), .msk_a0b2(din_2_msk_ab2), .msk_a0b3(din_2_msk_ab3),
           .msk_a0b0_1sc(din_2_msk_ab0_1sc), .msk_a0b1_1sc(din_2_msk_ab1_1sc), .msk_a0b2_1sc(din_2_msk_ab2_1sc), .msk_a0b3_1sc(din_2_msk_ab3_1sc),

           .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2),
           .a1b0_1sc(din_4_ab0_1sc), .a1b1_1sc(din_4_ab1_1sc), .a1b2_1sc(din_4_ab2_1sc),
           .msk_a1b0(din_4_msk_ab0), .msk_a1b1(din_4_msk_ab1), .msk_a1b2(din_4_msk_ab2),
           .msk_a1b0_1sc(din_4_msk_ab0_1sc), .msk_a1b1_1sc(din_4_msk_ab1_1sc), .msk_a1b2_1sc(din_4_msk_ab2_1sc),

           .a2b0(din_6_ab0), .a2b1(din_6_ab1),
           .a2b0_1sc(din_6_ab0_1sc), .a2b1_1sc(din_6_ab1_1sc),
           .msk_a2b0(din_6_msk_ab0), .msk_a2b1(din_6_msk_ab1),
           .msk_a2b0_1sc(din_6_msk_ab0_1sc), .msk_a2b1_1sc(din_6_msk_ab1_1sc),
           
           .a3b0(din_8_ab0),
           .a3b0_1sc(din_8_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_3_calc (
           .clk(clk), .sign(din_signs_reg[3]), 
           .p(addr_0_3),
           .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
           .a0b0_1sc(din_3_ab0_1sc), .a0b1_1sc(din_3_ab1_1sc), .a0b2_1sc(din_3_ab2_1sc), .a0b3_1sc(din_3_ab3_1sc),
           .msk_a0b0(din_3_msk_ab0), .msk_a0b1(din_3_msk_ab1), .msk_a0b2(din_3_msk_ab2), .msk_a0b3(din_3_msk_ab3),
           .msk_a0b0_1sc(din_3_msk_ab0_1sc), .msk_a0b1_1sc(din_3_msk_ab1_1sc), .msk_a0b2_1sc(din_3_msk_ab2_1sc), .msk_a0b3_1sc(din_3_msk_ab3_1sc),

           .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2),
           .a1b0_1sc(din_5_ab0_1sc), .a1b1_1sc(din_5_ab1_1sc), .a1b2_1sc(din_5_ab2_1sc),
           .msk_a1b0(din_5_msk_ab0), .msk_a1b1(din_5_msk_ab1), .msk_a1b2(din_5_msk_ab2),
           .msk_a1b0_1sc(din_5_msk_ab0_1sc), .msk_a1b1_1sc(din_5_msk_ab1_1sc), .msk_a1b2_1sc(din_5_msk_ab2_1sc),

           .a2b0(din_7_ab0), .a2b1(din_7_ab1),
           .a2b0_1sc(din_7_ab0_1sc), .a2b1_1sc(din_7_ab1_1sc),
           .msk_a2b0(din_7_msk_ab0), .msk_a2b1(din_7_msk_ab1),
           .msk_a2b0_1sc(din_7_msk_ab0_1sc), .msk_a2b1_1sc(din_7_msk_ab1_1sc),
           
           .a3b0(din_9_ab0),
           .a3b0_1sc(din_9_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_4_calc (
           .clk(clk), .sign(din_signs_reg[4]), 
           .p(addr_0_4),
           .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
           .a0b0_1sc(din_4_ab0_1sc), .a0b1_1sc(din_4_ab1_1sc), .a0b2_1sc(din_4_ab2_1sc), .a0b3_1sc(din_4_ab3_1sc),
           .msk_a0b0(din_4_msk_ab0), .msk_a0b1(din_4_msk_ab1), .msk_a0b2(din_4_msk_ab2), .msk_a0b3(din_4_msk_ab3),
           .msk_a0b0_1sc(din_4_msk_ab0_1sc), .msk_a0b1_1sc(din_4_msk_ab1_1sc), .msk_a0b2_1sc(din_4_msk_ab2_1sc), .msk_a0b3_1sc(din_4_msk_ab3_1sc),

           .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2),
           .a1b0_1sc(din_6_ab0_1sc), .a1b1_1sc(din_6_ab1_1sc), .a1b2_1sc(din_6_ab2_1sc),
           .msk_a1b0(din_6_msk_ab0), .msk_a1b1(din_6_msk_ab1), .msk_a1b2(din_6_msk_ab2),
           .msk_a1b0_1sc(din_6_msk_ab0_1sc), .msk_a1b1_1sc(din_6_msk_ab1_1sc), .msk_a1b2_1sc(din_6_msk_ab2_1sc),

           .a2b0(din_8_ab0), .a2b1(din_8_ab1),
           .a2b0_1sc(din_8_ab0_1sc), .a2b1_1sc(din_8_ab1_1sc),
           .msk_a2b0(din_8_msk_ab0), .msk_a2b1(din_8_msk_ab1),
           .msk_a2b0_1sc(din_8_msk_ab0_1sc), .msk_a2b1_1sc(din_8_msk_ab1_1sc),
           
           .a3b0(din_10_ab0),
           .a3b0_1sc(din_10_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_5_calc (
           .clk(clk), .sign(din_signs_reg[5]), 
           .p(addr_0_5),
           .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
           .a0b0_1sc(din_5_ab0_1sc), .a0b1_1sc(din_5_ab1_1sc), .a0b2_1sc(din_5_ab2_1sc), .a0b3_1sc(din_5_ab3_1sc),
           .msk_a0b0(din_5_msk_ab0), .msk_a0b1(din_5_msk_ab1), .msk_a0b2(din_5_msk_ab2), .msk_a0b3(din_5_msk_ab3),
           .msk_a0b0_1sc(din_5_msk_ab0_1sc), .msk_a0b1_1sc(din_5_msk_ab1_1sc), .msk_a0b2_1sc(din_5_msk_ab2_1sc), .msk_a0b3_1sc(din_5_msk_ab3_1sc),

           .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2),
           .a1b0_1sc(din_7_ab0_1sc), .a1b1_1sc(din_7_ab1_1sc), .a1b2_1sc(din_7_ab2_1sc),
           .msk_a1b0(din_7_msk_ab0), .msk_a1b1(din_7_msk_ab1), .msk_a1b2(din_7_msk_ab2),
           .msk_a1b0_1sc(din_7_msk_ab0_1sc), .msk_a1b1_1sc(din_7_msk_ab1_1sc), .msk_a1b2_1sc(din_7_msk_ab2_1sc),

           .a2b0(din_9_ab0), .a2b1(din_9_ab1),
           .a2b0_1sc(din_9_ab0_1sc), .a2b1_1sc(din_9_ab1_1sc),
           .msk_a2b0(din_9_msk_ab0), .msk_a2b1(din_9_msk_ab1),
           .msk_a2b0_1sc(din_9_msk_ab0_1sc), .msk_a2b1_1sc(din_9_msk_ab1_1sc),
           
           .a3b0(din_11_ab0),
           .a3b0_1sc(din_11_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_6_calc (
           .clk(clk), .sign(din_signs_reg[6]), 
           .p(addr_0_6),
           .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
           .a0b0_1sc(din_6_ab0_1sc), .a0b1_1sc(din_6_ab1_1sc), .a0b2_1sc(din_6_ab2_1sc), .a0b3_1sc(din_6_ab3_1sc),
           .msk_a0b0(din_6_msk_ab0), .msk_a0b1(din_6_msk_ab1), .msk_a0b2(din_6_msk_ab2), .msk_a0b3(din_6_msk_ab3),
           .msk_a0b0_1sc(din_6_msk_ab0_1sc), .msk_a0b1_1sc(din_6_msk_ab1_1sc), .msk_a0b2_1sc(din_6_msk_ab2_1sc), .msk_a0b3_1sc(din_6_msk_ab3_1sc),

           .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2),
           .a1b0_1sc(din_8_ab0_1sc), .a1b1_1sc(din_8_ab1_1sc), .a1b2_1sc(din_8_ab2_1sc),
           .msk_a1b0(din_8_msk_ab0), .msk_a1b1(din_8_msk_ab1), .msk_a1b2(din_8_msk_ab2),
           .msk_a1b0_1sc(din_8_msk_ab0_1sc), .msk_a1b1_1sc(din_8_msk_ab1_1sc), .msk_a1b2_1sc(din_8_msk_ab2_1sc),

           .a2b0(din_10_ab0), .a2b1(din_10_ab1),
           .a2b0_1sc(din_10_ab0_1sc), .a2b1_1sc(din_10_ab1_1sc),
           .msk_a2b0(din_10_msk_ab0), .msk_a2b1(din_10_msk_ab1),
           .msk_a2b0_1sc(din_10_msk_ab0_1sc), .msk_a2b1_1sc(din_10_msk_ab1_1sc),
           
           .a3b0(din_12_ab0),
           .a3b0_1sc(din_12_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_7_calc (
           .clk(clk), .sign(din_signs_reg[7]), 
           .p(addr_0_7),
           .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
           .a0b0_1sc(din_7_ab0_1sc), .a0b1_1sc(din_7_ab1_1sc), .a0b2_1sc(din_7_ab2_1sc), .a0b3_1sc(din_7_ab3_1sc),
           .msk_a0b0(din_7_msk_ab0), .msk_a0b1(din_7_msk_ab1), .msk_a0b2(din_7_msk_ab2), .msk_a0b3(din_7_msk_ab3),
           .msk_a0b0_1sc(din_7_msk_ab0_1sc), .msk_a0b1_1sc(din_7_msk_ab1_1sc), .msk_a0b2_1sc(din_7_msk_ab2_1sc), .msk_a0b3_1sc(din_7_msk_ab3_1sc),

           .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2),
           .a1b0_1sc(din_9_ab0_1sc), .a1b1_1sc(din_9_ab1_1sc), .a1b2_1sc(din_9_ab2_1sc),
           .msk_a1b0(din_9_msk_ab0), .msk_a1b1(din_9_msk_ab1), .msk_a1b2(din_9_msk_ab2),
           .msk_a1b0_1sc(din_9_msk_ab0_1sc), .msk_a1b1_1sc(din_9_msk_ab1_1sc), .msk_a1b2_1sc(din_9_msk_ab2_1sc),

           .a2b0(din_11_ab0), .a2b1(din_11_ab1),
           .a2b0_1sc(din_11_ab0_1sc), .a2b1_1sc(din_11_ab1_1sc),
           .msk_a2b0(din_11_msk_ab0), .msk_a2b1(din_11_msk_ab1),
           .msk_a2b0_1sc(din_11_msk_ab0_1sc), .msk_a2b1_1sc(din_11_msk_ab1_1sc),
           
           .a3b0(din_13_ab0),
           .a3b0_1sc(din_13_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_8_calc (
           .clk(clk), .sign(din_signs_reg[8]), 
           .p(addr_0_8),
           .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
           .a0b0_1sc(din_8_ab0_1sc), .a0b1_1sc(din_8_ab1_1sc), .a0b2_1sc(din_8_ab2_1sc), .a0b3_1sc(din_8_ab3_1sc),
           .msk_a0b0(din_8_msk_ab0), .msk_a0b1(din_8_msk_ab1), .msk_a0b2(din_8_msk_ab2), .msk_a0b3(din_8_msk_ab3),
           .msk_a0b0_1sc(din_8_msk_ab0_1sc), .msk_a0b1_1sc(din_8_msk_ab1_1sc), .msk_a0b2_1sc(din_8_msk_ab2_1sc), .msk_a0b3_1sc(din_8_msk_ab3_1sc),

           .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2),
           .a1b0_1sc(din_10_ab0_1sc), .a1b1_1sc(din_10_ab1_1sc), .a1b2_1sc(din_10_ab2_1sc),
           .msk_a1b0(din_10_msk_ab0), .msk_a1b1(din_10_msk_ab1), .msk_a1b2(din_10_msk_ab2),
           .msk_a1b0_1sc(din_10_msk_ab0_1sc), .msk_a1b1_1sc(din_10_msk_ab1_1sc), .msk_a1b2_1sc(din_10_msk_ab2_1sc),

           .a2b0(din_12_ab0), .a2b1(din_12_ab1),
           .a2b0_1sc(din_12_ab0_1sc), .a2b1_1sc(din_12_ab1_1sc),
           .msk_a2b0(din_12_msk_ab0), .msk_a2b1(din_12_msk_ab1),
           .msk_a2b0_1sc(din_12_msk_ab0_1sc), .msk_a2b1_1sc(din_12_msk_ab1_1sc),
           
           .a3b0(din_14_ab0),
           .a3b0_1sc(din_14_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_9_calc (
           .clk(clk), .sign(din_signs_reg[9]), 
           .p(addr_0_9),
           .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
           .a0b0_1sc(din_9_ab0_1sc), .a0b1_1sc(din_9_ab1_1sc), .a0b2_1sc(din_9_ab2_1sc), .a0b3_1sc(din_9_ab3_1sc),
           .msk_a0b0(din_9_msk_ab0), .msk_a0b1(din_9_msk_ab1), .msk_a0b2(din_9_msk_ab2), .msk_a0b3(din_9_msk_ab3),
           .msk_a0b0_1sc(din_9_msk_ab0_1sc), .msk_a0b1_1sc(din_9_msk_ab1_1sc), .msk_a0b2_1sc(din_9_msk_ab2_1sc), .msk_a0b3_1sc(din_9_msk_ab3_1sc),

           .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2),
           .a1b0_1sc(din_11_ab0_1sc), .a1b1_1sc(din_11_ab1_1sc), .a1b2_1sc(din_11_ab2_1sc),
           .msk_a1b0(din_11_msk_ab0), .msk_a1b1(din_11_msk_ab1), .msk_a1b2(din_11_msk_ab2),
           .msk_a1b0_1sc(din_11_msk_ab0_1sc), .msk_a1b1_1sc(din_11_msk_ab1_1sc), .msk_a1b2_1sc(din_11_msk_ab2_1sc),

           .a2b0(din_13_ab0), .a2b1(din_13_ab1),
           .a2b0_1sc(din_13_ab0_1sc), .a2b1_1sc(din_13_ab1_1sc),
           .msk_a2b0(din_13_msk_ab0), .msk_a2b1(din_13_msk_ab1),
           .msk_a2b0_1sc(din_13_msk_ab0_1sc), .msk_a2b1_1sc(din_13_msk_ab1_1sc),
           
           .a3b0(din_15_ab0),
           .a3b0_1sc(din_15_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_10_calc (
           .clk(clk), .sign(din_signs_reg[10]), 
           .p(addr_0_10),
           .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
           .a0b0_1sc(din_10_ab0_1sc), .a0b1_1sc(din_10_ab1_1sc), .a0b2_1sc(din_10_ab2_1sc), .a0b3_1sc(din_10_ab3_1sc),
           .msk_a0b0(din_10_msk_ab0), .msk_a0b1(din_10_msk_ab1), .msk_a0b2(din_10_msk_ab2), .msk_a0b3(din_10_msk_ab3),
           .msk_a0b0_1sc(din_10_msk_ab0_1sc), .msk_a0b1_1sc(din_10_msk_ab1_1sc), .msk_a0b2_1sc(din_10_msk_ab2_1sc), .msk_a0b3_1sc(din_10_msk_ab3_1sc),

           .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2),
           .a1b0_1sc(din_12_ab0_1sc), .a1b1_1sc(din_12_ab1_1sc), .a1b2_1sc(din_12_ab2_1sc),
           .msk_a1b0(din_12_msk_ab0), .msk_a1b1(din_12_msk_ab1), .msk_a1b2(din_12_msk_ab2),
           .msk_a1b0_1sc(din_12_msk_ab0_1sc), .msk_a1b1_1sc(din_12_msk_ab1_1sc), .msk_a1b2_1sc(din_12_msk_ab2_1sc),

           .a2b0(din_14_ab0), .a2b1(din_14_ab1),
           .a2b0_1sc(din_14_ab0_1sc), .a2b1_1sc(din_14_ab1_1sc),
           .msk_a2b0(din_14_msk_ab0), .msk_a2b1(din_14_msk_ab1),
           .msk_a2b0_1sc(din_14_msk_ab0_1sc), .msk_a2b1_1sc(din_14_msk_ab1_1sc),
           
           .a3b0(din_16_ab0),
           .a3b0_1sc(din_16_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_11_calc (
           .clk(clk), .sign(din_signs_reg[11]), 
           .p(addr_0_11),
           .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
           .a0b0_1sc(din_11_ab0_1sc), .a0b1_1sc(din_11_ab1_1sc), .a0b2_1sc(din_11_ab2_1sc), .a0b3_1sc(din_11_ab3_1sc),
           .msk_a0b0(din_11_msk_ab0), .msk_a0b1(din_11_msk_ab1), .msk_a0b2(din_11_msk_ab2), .msk_a0b3(din_11_msk_ab3),
           .msk_a0b0_1sc(din_11_msk_ab0_1sc), .msk_a0b1_1sc(din_11_msk_ab1_1sc), .msk_a0b2_1sc(din_11_msk_ab2_1sc), .msk_a0b3_1sc(din_11_msk_ab3_1sc),

           .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2),
           .a1b0_1sc(din_13_ab0_1sc), .a1b1_1sc(din_13_ab1_1sc), .a1b2_1sc(din_13_ab2_1sc),
           .msk_a1b0(din_13_msk_ab0), .msk_a1b1(din_13_msk_ab1), .msk_a1b2(din_13_msk_ab2),
           .msk_a1b0_1sc(din_13_msk_ab0_1sc), .msk_a1b1_1sc(din_13_msk_ab1_1sc), .msk_a1b2_1sc(din_13_msk_ab2_1sc),

           .a2b0(din_15_ab0), .a2b1(din_15_ab1),
           .a2b0_1sc(din_15_ab0_1sc), .a2b1_1sc(din_15_ab1_1sc),
           .msk_a2b0(din_15_msk_ab0), .msk_a2b1(din_15_msk_ab1),
           .msk_a2b0_1sc(din_15_msk_ab0_1sc), .msk_a2b1_1sc(din_15_msk_ab1_1sc),
           
           .a3b0(din_17_ab0),
           .a3b0_1sc(din_17_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_12_calc (
           .clk(clk), .sign(din_signs_reg[12]), 
           .p(addr_0_12),
           .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
           .a0b0_1sc(din_12_ab0_1sc), .a0b1_1sc(din_12_ab1_1sc), .a0b2_1sc(din_12_ab2_1sc), .a0b3_1sc(din_12_ab3_1sc),
           .msk_a0b0(din_12_msk_ab0), .msk_a0b1(din_12_msk_ab1), .msk_a0b2(din_12_msk_ab2), .msk_a0b3(din_12_msk_ab3),
           .msk_a0b0_1sc(din_12_msk_ab0_1sc), .msk_a0b1_1sc(din_12_msk_ab1_1sc), .msk_a0b2_1sc(din_12_msk_ab2_1sc), .msk_a0b3_1sc(din_12_msk_ab3_1sc),

           .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2),
           .a1b0_1sc(din_14_ab0_1sc), .a1b1_1sc(din_14_ab1_1sc), .a1b2_1sc(din_14_ab2_1sc),
           .msk_a1b0(din_14_msk_ab0), .msk_a1b1(din_14_msk_ab1), .msk_a1b2(din_14_msk_ab2),
           .msk_a1b0_1sc(din_14_msk_ab0_1sc), .msk_a1b1_1sc(din_14_msk_ab1_1sc), .msk_a1b2_1sc(din_14_msk_ab2_1sc),

           .a2b0(din_16_ab0), .a2b1(din_16_ab1),
           .a2b0_1sc(din_16_ab0_1sc), .a2b1_1sc(din_16_ab1_1sc),
           .msk_a2b0(din_16_msk_ab0), .msk_a2b1(din_16_msk_ab1),
           .msk_a2b0_1sc(din_16_msk_ab0_1sc), .msk_a2b1_1sc(din_16_msk_ab1_1sc),
           
           .a3b0(din_18_ab0),
           .a3b0_1sc(din_18_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_13_calc (
           .clk(clk), .sign(din_signs_reg[13]), 
           .p(addr_0_13),
           .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
           .a0b0_1sc(din_13_ab0_1sc), .a0b1_1sc(din_13_ab1_1sc), .a0b2_1sc(din_13_ab2_1sc), .a0b3_1sc(din_13_ab3_1sc),
           .msk_a0b0(din_13_msk_ab0), .msk_a0b1(din_13_msk_ab1), .msk_a0b2(din_13_msk_ab2), .msk_a0b3(din_13_msk_ab3),
           .msk_a0b0_1sc(din_13_msk_ab0_1sc), .msk_a0b1_1sc(din_13_msk_ab1_1sc), .msk_a0b2_1sc(din_13_msk_ab2_1sc), .msk_a0b3_1sc(din_13_msk_ab3_1sc),

           .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2),
           .a1b0_1sc(din_15_ab0_1sc), .a1b1_1sc(din_15_ab1_1sc), .a1b2_1sc(din_15_ab2_1sc),
           .msk_a1b0(din_15_msk_ab0), .msk_a1b1(din_15_msk_ab1), .msk_a1b2(din_15_msk_ab2),
           .msk_a1b0_1sc(din_15_msk_ab0_1sc), .msk_a1b1_1sc(din_15_msk_ab1_1sc), .msk_a1b2_1sc(din_15_msk_ab2_1sc),

           .a2b0(din_17_ab0), .a2b1(din_17_ab1),
           .a2b0_1sc(din_17_ab0_1sc), .a2b1_1sc(din_17_ab1_1sc),
           .msk_a2b0(din_17_msk_ab0), .msk_a2b1(din_17_msk_ab1),
           .msk_a2b0_1sc(din_17_msk_ab0_1sc), .msk_a2b1_1sc(din_17_msk_ab1_1sc),
           
           .a3b0(din_19_ab0),
           .a3b0_1sc(din_19_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_14_calc (
           .clk(clk), .sign(din_signs_reg[14]), 
           .p(addr_0_14),
           .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
           .a0b0_1sc(din_14_ab0_1sc), .a0b1_1sc(din_14_ab1_1sc), .a0b2_1sc(din_14_ab2_1sc), .a0b3_1sc(din_14_ab3_1sc),
           .msk_a0b0(din_14_msk_ab0), .msk_a0b1(din_14_msk_ab1), .msk_a0b2(din_14_msk_ab2), .msk_a0b3(din_14_msk_ab3),
           .msk_a0b0_1sc(din_14_msk_ab0_1sc), .msk_a0b1_1sc(din_14_msk_ab1_1sc), .msk_a0b2_1sc(din_14_msk_ab2_1sc), .msk_a0b3_1sc(din_14_msk_ab3_1sc),

           .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2),
           .a1b0_1sc(din_16_ab0_1sc), .a1b1_1sc(din_16_ab1_1sc), .a1b2_1sc(din_16_ab2_1sc),
           .msk_a1b0(din_16_msk_ab0), .msk_a1b1(din_16_msk_ab1), .msk_a1b2(din_16_msk_ab2),
           .msk_a1b0_1sc(din_16_msk_ab0_1sc), .msk_a1b1_1sc(din_16_msk_ab1_1sc), .msk_a1b2_1sc(din_16_msk_ab2_1sc),

           .a2b0(din_18_ab0), .a2b1(din_18_ab1),
           .a2b0_1sc(din_18_ab0_1sc), .a2b1_1sc(din_18_ab1_1sc),
           .msk_a2b0(din_18_msk_ab0), .msk_a2b1(din_18_msk_ab1),
           .msk_a2b0_1sc(din_18_msk_ab0_1sc), .msk_a2b1_1sc(din_18_msk_ab1_1sc),
           
           .a3b0(din_20_ab0),
           .a3b0_1sc(din_20_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_15_calc (
           .clk(clk), .sign(din_signs_reg[15]), 
           .p(addr_0_15),
           .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
           .a0b0_1sc(din_15_ab0_1sc), .a0b1_1sc(din_15_ab1_1sc), .a0b2_1sc(din_15_ab2_1sc), .a0b3_1sc(din_15_ab3_1sc),
           .msk_a0b0(din_15_msk_ab0), .msk_a0b1(din_15_msk_ab1), .msk_a0b2(din_15_msk_ab2), .msk_a0b3(din_15_msk_ab3),
           .msk_a0b0_1sc(din_15_msk_ab0_1sc), .msk_a0b1_1sc(din_15_msk_ab1_1sc), .msk_a0b2_1sc(din_15_msk_ab2_1sc), .msk_a0b3_1sc(din_15_msk_ab3_1sc),

           .a1b0(din_17_ab0), .a1b1(din_17_ab1), .a1b2(din_17_ab2),
           .a1b0_1sc(din_17_ab0_1sc), .a1b1_1sc(din_17_ab1_1sc), .a1b2_1sc(din_17_ab2_1sc),
           .msk_a1b0(din_17_msk_ab0), .msk_a1b1(din_17_msk_ab1), .msk_a1b2(din_17_msk_ab2),
           .msk_a1b0_1sc(din_17_msk_ab0_1sc), .msk_a1b1_1sc(din_17_msk_ab1_1sc), .msk_a1b2_1sc(din_17_msk_ab2_1sc),

           .a2b0(din_19_ab0), .a2b1(din_19_ab1),
           .a2b0_1sc(din_19_ab0_1sc), .a2b1_1sc(din_19_ab1_1sc),
           .msk_a2b0(din_19_msk_ab0), .msk_a2b1(din_19_msk_ab1),
           .msk_a2b0_1sc(din_19_msk_ab0_1sc), .msk_a2b1_1sc(din_19_msk_ab1_1sc),
           
           .a3b0(din_21_ab0),
           .a3b0_1sc(din_21_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_16_calc (
           .clk(clk), .sign(din_signs_reg[16]), 
           .p(addr_0_16),
           .a0b0(din_16_ab0), .a0b1(din_16_ab1), .a0b2(din_16_ab2), .a0b3(din_16_ab3),
           .a0b0_1sc(din_16_ab0_1sc), .a0b1_1sc(din_16_ab1_1sc), .a0b2_1sc(din_16_ab2_1sc), .a0b3_1sc(din_16_ab3_1sc),
           .msk_a0b0(din_16_msk_ab0), .msk_a0b1(din_16_msk_ab1), .msk_a0b2(din_16_msk_ab2), .msk_a0b3(din_16_msk_ab3),
           .msk_a0b0_1sc(din_16_msk_ab0_1sc), .msk_a0b1_1sc(din_16_msk_ab1_1sc), .msk_a0b2_1sc(din_16_msk_ab2_1sc), .msk_a0b3_1sc(din_16_msk_ab3_1sc),

           .a1b0(din_18_ab0), .a1b1(din_18_ab1), .a1b2(din_18_ab2),
           .a1b0_1sc(din_18_ab0_1sc), .a1b1_1sc(din_18_ab1_1sc), .a1b2_1sc(din_18_ab2_1sc),
           .msk_a1b0(din_18_msk_ab0), .msk_a1b1(din_18_msk_ab1), .msk_a1b2(din_18_msk_ab2),
           .msk_a1b0_1sc(din_18_msk_ab0_1sc), .msk_a1b1_1sc(din_18_msk_ab1_1sc), .msk_a1b2_1sc(din_18_msk_ab2_1sc),

           .a2b0(din_20_ab0), .a2b1(din_20_ab1),
           .a2b0_1sc(din_20_ab0_1sc), .a2b1_1sc(din_20_ab1_1sc),
           .msk_a2b0(din_20_msk_ab0), .msk_a2b1(din_20_msk_ab1),
           .msk_a2b0_1sc(din_20_msk_ab0_1sc), .msk_a2b1_1sc(din_20_msk_ab1_1sc),
           
           .a3b0(din_22_ab0),
           .a3b0_1sc(din_22_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_17_calc (
           .clk(clk), .sign(din_signs_reg[17]), 
           .p(addr_0_17),
           .a0b0(din_17_ab0), .a0b1(din_17_ab1), .a0b2(din_17_ab2), .a0b3(din_17_ab3),
           .a0b0_1sc(din_17_ab0_1sc), .a0b1_1sc(din_17_ab1_1sc), .a0b2_1sc(din_17_ab2_1sc), .a0b3_1sc(din_17_ab3_1sc),
           .msk_a0b0(din_17_msk_ab0), .msk_a0b1(din_17_msk_ab1), .msk_a0b2(din_17_msk_ab2), .msk_a0b3(din_17_msk_ab3),
           .msk_a0b0_1sc(din_17_msk_ab0_1sc), .msk_a0b1_1sc(din_17_msk_ab1_1sc), .msk_a0b2_1sc(din_17_msk_ab2_1sc), .msk_a0b3_1sc(din_17_msk_ab3_1sc),

           .a1b0(din_19_ab0), .a1b1(din_19_ab1), .a1b2(din_19_ab2),
           .a1b0_1sc(din_19_ab0_1sc), .a1b1_1sc(din_19_ab1_1sc), .a1b2_1sc(din_19_ab2_1sc),
           .msk_a1b0(din_19_msk_ab0), .msk_a1b1(din_19_msk_ab1), .msk_a1b2(din_19_msk_ab2),
           .msk_a1b0_1sc(din_19_msk_ab0_1sc), .msk_a1b1_1sc(din_19_msk_ab1_1sc), .msk_a1b2_1sc(din_19_msk_ab2_1sc),

           .a2b0(din_21_ab0), .a2b1(din_21_ab1),
           .a2b0_1sc(din_21_ab0_1sc), .a2b1_1sc(din_21_ab1_1sc),
           .msk_a2b0(din_21_msk_ab0), .msk_a2b1(din_21_msk_ab1),
           .msk_a2b0_1sc(din_21_msk_ab0_1sc), .msk_a2b1_1sc(din_21_msk_ab1_1sc),
           
           .a3b0(din_23_ab0),
           .a3b0_1sc(din_23_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_18_calc (
           .clk(clk), .sign(din_signs_reg[18]), 
           .p(addr_0_18),
           .a0b0(din_18_ab0), .a0b1(din_18_ab1), .a0b2(din_18_ab2), .a0b3(din_18_ab3),
           .a0b0_1sc(din_18_ab0_1sc), .a0b1_1sc(din_18_ab1_1sc), .a0b2_1sc(din_18_ab2_1sc), .a0b3_1sc(din_18_ab3_1sc),
           .msk_a0b0(din_18_msk_ab0), .msk_a0b1(din_18_msk_ab1), .msk_a0b2(din_18_msk_ab2), .msk_a0b3(din_18_msk_ab3),
           .msk_a0b0_1sc(din_18_msk_ab0_1sc), .msk_a0b1_1sc(din_18_msk_ab1_1sc), .msk_a0b2_1sc(din_18_msk_ab2_1sc), .msk_a0b3_1sc(din_18_msk_ab3_1sc),

           .a1b0(din_20_ab0), .a1b1(din_20_ab1), .a1b2(din_20_ab2),
           .a1b0_1sc(din_20_ab0_1sc), .a1b1_1sc(din_20_ab1_1sc), .a1b2_1sc(din_20_ab2_1sc),
           .msk_a1b0(din_20_msk_ab0), .msk_a1b1(din_20_msk_ab1), .msk_a1b2(din_20_msk_ab2),
           .msk_a1b0_1sc(din_20_msk_ab0_1sc), .msk_a1b1_1sc(din_20_msk_ab1_1sc), .msk_a1b2_1sc(din_20_msk_ab2_1sc),

           .a2b0(din_22_ab0), .a2b1(din_22_ab1),
           .a2b0_1sc(din_22_ab0_1sc), .a2b1_1sc(din_22_ab1_1sc),
           .msk_a2b0(din_22_msk_ab0), .msk_a2b1(din_22_msk_ab1),
           .msk_a2b0_1sc(din_22_msk_ab0_1sc), .msk_a2b1_1sc(din_22_msk_ab1_1sc),
           
           .a3b0(din_24_ab0),
           .a3b0_1sc(din_24_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_19_calc (
           .clk(clk), .sign(din_signs_reg[19]), 
           .p(addr_0_19),
           .a0b0(din_19_ab0), .a0b1(din_19_ab1), .a0b2(din_19_ab2), .a0b3(din_19_ab3),
           .a0b0_1sc(din_19_ab0_1sc), .a0b1_1sc(din_19_ab1_1sc), .a0b2_1sc(din_19_ab2_1sc), .a0b3_1sc(din_19_ab3_1sc),
           .msk_a0b0(din_19_msk_ab0), .msk_a0b1(din_19_msk_ab1), .msk_a0b2(din_19_msk_ab2), .msk_a0b3(din_19_msk_ab3),
           .msk_a0b0_1sc(din_19_msk_ab0_1sc), .msk_a0b1_1sc(din_19_msk_ab1_1sc), .msk_a0b2_1sc(din_19_msk_ab2_1sc), .msk_a0b3_1sc(din_19_msk_ab3_1sc),

           .a1b0(din_21_ab0), .a1b1(din_21_ab1), .a1b2(din_21_ab2),
           .a1b0_1sc(din_21_ab0_1sc), .a1b1_1sc(din_21_ab1_1sc), .a1b2_1sc(din_21_ab2_1sc),
           .msk_a1b0(din_21_msk_ab0), .msk_a1b1(din_21_msk_ab1), .msk_a1b2(din_21_msk_ab2),
           .msk_a1b0_1sc(din_21_msk_ab0_1sc), .msk_a1b1_1sc(din_21_msk_ab1_1sc), .msk_a1b2_1sc(din_21_msk_ab2_1sc),

           .a2b0(din_23_ab0), .a2b1(din_23_ab1),
           .a2b0_1sc(din_23_ab0_1sc), .a2b1_1sc(din_23_ab1_1sc),
           .msk_a2b0(din_23_msk_ab0), .msk_a2b1(din_23_msk_ab1),
           .msk_a2b0_1sc(din_23_msk_ab0_1sc), .msk_a2b1_1sc(din_23_msk_ab1_1sc),
           
           .a3b0(din_25_ab0),
           .a3b0_1sc(din_25_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_20_calc (
           .clk(clk), .sign(din_signs_reg[20]), 
           .p(addr_0_20),
           .a0b0(din_20_ab0), .a0b1(din_20_ab1), .a0b2(din_20_ab2), .a0b3(din_20_ab3),
           .a0b0_1sc(din_20_ab0_1sc), .a0b1_1sc(din_20_ab1_1sc), .a0b2_1sc(din_20_ab2_1sc), .a0b3_1sc(din_20_ab3_1sc),
           .msk_a0b0(din_20_msk_ab0), .msk_a0b1(din_20_msk_ab1), .msk_a0b2(din_20_msk_ab2), .msk_a0b3(din_20_msk_ab3),
           .msk_a0b0_1sc(din_20_msk_ab0_1sc), .msk_a0b1_1sc(din_20_msk_ab1_1sc), .msk_a0b2_1sc(din_20_msk_ab2_1sc), .msk_a0b3_1sc(din_20_msk_ab3_1sc),

           .a1b0(din_22_ab0), .a1b1(din_22_ab1), .a1b2(din_22_ab2),
           .a1b0_1sc(din_22_ab0_1sc), .a1b1_1sc(din_22_ab1_1sc), .a1b2_1sc(din_22_ab2_1sc),
           .msk_a1b0(din_22_msk_ab0), .msk_a1b1(din_22_msk_ab1), .msk_a1b2(din_22_msk_ab2),
           .msk_a1b0_1sc(din_22_msk_ab0_1sc), .msk_a1b1_1sc(din_22_msk_ab1_1sc), .msk_a1b2_1sc(din_22_msk_ab2_1sc),

           .a2b0(din_24_ab0), .a2b1(din_24_ab1),
           .a2b0_1sc(din_24_ab0_1sc), .a2b1_1sc(din_24_ab1_1sc),
           .msk_a2b0(din_24_msk_ab0), .msk_a2b1(din_24_msk_ab1),
           .msk_a2b0_1sc(din_24_msk_ab0_1sc), .msk_a2b1_1sc(din_24_msk_ab1_1sc),
           
           .a3b0(din_26_ab0),
           .a3b0_1sc(din_26_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_21_calc (
           .clk(clk), .sign(din_signs_reg[21]), 
           .p(addr_0_21),
           .a0b0(din_21_ab0), .a0b1(din_21_ab1), .a0b2(din_21_ab2), .a0b3(din_21_ab3),
           .a0b0_1sc(din_21_ab0_1sc), .a0b1_1sc(din_21_ab1_1sc), .a0b2_1sc(din_21_ab2_1sc), .a0b3_1sc(din_21_ab3_1sc),
           .msk_a0b0(din_21_msk_ab0), .msk_a0b1(din_21_msk_ab1), .msk_a0b2(din_21_msk_ab2), .msk_a0b3(din_21_msk_ab3),
           .msk_a0b0_1sc(din_21_msk_ab0_1sc), .msk_a0b1_1sc(din_21_msk_ab1_1sc), .msk_a0b2_1sc(din_21_msk_ab2_1sc), .msk_a0b3_1sc(din_21_msk_ab3_1sc),

           .a1b0(din_23_ab0), .a1b1(din_23_ab1), .a1b2(din_23_ab2),
           .a1b0_1sc(din_23_ab0_1sc), .a1b1_1sc(din_23_ab1_1sc), .a1b2_1sc(din_23_ab2_1sc),
           .msk_a1b0(din_23_msk_ab0), .msk_a1b1(din_23_msk_ab1), .msk_a1b2(din_23_msk_ab2),
           .msk_a1b0_1sc(din_23_msk_ab0_1sc), .msk_a1b1_1sc(din_23_msk_ab1_1sc), .msk_a1b2_1sc(din_23_msk_ab2_1sc),

           .a2b0(din_25_ab0), .a2b1(din_25_ab1),
           .a2b0_1sc(din_25_ab0_1sc), .a2b1_1sc(din_25_ab1_1sc),
           .msk_a2b0(din_25_msk_ab0), .msk_a2b1(din_25_msk_ab1),
           .msk_a2b0_1sc(din_25_msk_ab0_1sc), .msk_a2b1_1sc(din_25_msk_ab1_1sc),
           
           .a3b0(din_27_ab0),
           .a3b0_1sc(din_27_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_22_calc (
           .clk(clk), .sign(din_signs_reg[22]), 
           .p(addr_0_22),
           .a0b0(din_22_ab0), .a0b1(din_22_ab1), .a0b2(din_22_ab2), .a0b3(din_22_ab3),
           .a0b0_1sc(din_22_ab0_1sc), .a0b1_1sc(din_22_ab1_1sc), .a0b2_1sc(din_22_ab2_1sc), .a0b3_1sc(din_22_ab3_1sc),
           .msk_a0b0(din_22_msk_ab0), .msk_a0b1(din_22_msk_ab1), .msk_a0b2(din_22_msk_ab2), .msk_a0b3(din_22_msk_ab3),
           .msk_a0b0_1sc(din_22_msk_ab0_1sc), .msk_a0b1_1sc(din_22_msk_ab1_1sc), .msk_a0b2_1sc(din_22_msk_ab2_1sc), .msk_a0b3_1sc(din_22_msk_ab3_1sc),

           .a1b0(din_24_ab0), .a1b1(din_24_ab1), .a1b2(din_24_ab2),
           .a1b0_1sc(din_24_ab0_1sc), .a1b1_1sc(din_24_ab1_1sc), .a1b2_1sc(din_24_ab2_1sc),
           .msk_a1b0(din_24_msk_ab0), .msk_a1b1(din_24_msk_ab1), .msk_a1b2(din_24_msk_ab2),
           .msk_a1b0_1sc(din_24_msk_ab0_1sc), .msk_a1b1_1sc(din_24_msk_ab1_1sc), .msk_a1b2_1sc(din_24_msk_ab2_1sc),

           .a2b0(din_26_ab0), .a2b1(din_26_ab1),
           .a2b0_1sc(din_26_ab0_1sc), .a2b1_1sc(din_26_ab1_1sc),
           .msk_a2b0(din_26_msk_ab0), .msk_a2b1(din_26_msk_ab1),
           .msk_a2b0_1sc(din_26_msk_ab0_1sc), .msk_a2b1_1sc(din_26_msk_ab1_1sc),
           
           .a3b0(din_28_ab0),
           .a3b0_1sc(din_28_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_23_calc (
           .clk(clk), .sign(din_signs_reg[23]), 
           .p(addr_0_23),
           .a0b0(din_23_ab0), .a0b1(din_23_ab1), .a0b2(din_23_ab2), .a0b3(din_23_ab3),
           .a0b0_1sc(din_23_ab0_1sc), .a0b1_1sc(din_23_ab1_1sc), .a0b2_1sc(din_23_ab2_1sc), .a0b3_1sc(din_23_ab3_1sc),
           .msk_a0b0(din_23_msk_ab0), .msk_a0b1(din_23_msk_ab1), .msk_a0b2(din_23_msk_ab2), .msk_a0b3(din_23_msk_ab3),
           .msk_a0b0_1sc(din_23_msk_ab0_1sc), .msk_a0b1_1sc(din_23_msk_ab1_1sc), .msk_a0b2_1sc(din_23_msk_ab2_1sc), .msk_a0b3_1sc(din_23_msk_ab3_1sc),

           .a1b0(din_25_ab0), .a1b1(din_25_ab1), .a1b2(din_25_ab2),
           .a1b0_1sc(din_25_ab0_1sc), .a1b1_1sc(din_25_ab1_1sc), .a1b2_1sc(din_25_ab2_1sc),
           .msk_a1b0(din_25_msk_ab0), .msk_a1b1(din_25_msk_ab1), .msk_a1b2(din_25_msk_ab2),
           .msk_a1b0_1sc(din_25_msk_ab0_1sc), .msk_a1b1_1sc(din_25_msk_ab1_1sc), .msk_a1b2_1sc(din_25_msk_ab2_1sc),

           .a2b0(din_27_ab0), .a2b1(din_27_ab1),
           .a2b0_1sc(din_27_ab0_1sc), .a2b1_1sc(din_27_ab1_1sc),
           .msk_a2b0(din_27_msk_ab0), .msk_a2b1(din_27_msk_ab1),
           .msk_a2b0_1sc(din_27_msk_ab0_1sc), .msk_a2b1_1sc(din_27_msk_ab1_1sc),
           
           .a3b0(din_29_ab0),
           .a3b0_1sc(din_29_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_24_calc (
           .clk(clk), .sign(din_signs_reg[24]), 
           .p(addr_0_24),
           .a0b0(din_24_ab0), .a0b1(din_24_ab1), .a0b2(din_24_ab2), .a0b3(din_24_ab3),
           .a0b0_1sc(din_24_ab0_1sc), .a0b1_1sc(din_24_ab1_1sc), .a0b2_1sc(din_24_ab2_1sc), .a0b3_1sc(din_24_ab3_1sc),
           .msk_a0b0(din_24_msk_ab0), .msk_a0b1(din_24_msk_ab1), .msk_a0b2(din_24_msk_ab2), .msk_a0b3(din_24_msk_ab3),
           .msk_a0b0_1sc(din_24_msk_ab0_1sc), .msk_a0b1_1sc(din_24_msk_ab1_1sc), .msk_a0b2_1sc(din_24_msk_ab2_1sc), .msk_a0b3_1sc(din_24_msk_ab3_1sc),

           .a1b0(din_26_ab0), .a1b1(din_26_ab1), .a1b2(din_26_ab2),
           .a1b0_1sc(din_26_ab0_1sc), .a1b1_1sc(din_26_ab1_1sc), .a1b2_1sc(din_26_ab2_1sc),
           .msk_a1b0(din_26_msk_ab0), .msk_a1b1(din_26_msk_ab1), .msk_a1b2(din_26_msk_ab2),
           .msk_a1b0_1sc(din_26_msk_ab0_1sc), .msk_a1b1_1sc(din_26_msk_ab1_1sc), .msk_a1b2_1sc(din_26_msk_ab2_1sc),

           .a2b0(din_28_ab0), .a2b1(din_28_ab1),
           .a2b0_1sc(din_28_ab0_1sc), .a2b1_1sc(din_28_ab1_1sc),
           .msk_a2b0(din_28_msk_ab0), .msk_a2b1(din_28_msk_ab1),
           .msk_a2b0_1sc(din_28_msk_ab0_1sc), .msk_a2b1_1sc(din_28_msk_ab1_1sc),
           
           .a3b0(din_30_ab0),
           .a3b0_1sc(din_30_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_25_calc (
           .clk(clk), .sign(din_signs_reg[25]), 
           .p(addr_0_25),
           .a0b0(din_25_ab0), .a0b1(din_25_ab1), .a0b2(din_25_ab2), .a0b3(din_25_ab3),
           .a0b0_1sc(din_25_ab0_1sc), .a0b1_1sc(din_25_ab1_1sc), .a0b2_1sc(din_25_ab2_1sc), .a0b3_1sc(din_25_ab3_1sc),
           .msk_a0b0(din_25_msk_ab0), .msk_a0b1(din_25_msk_ab1), .msk_a0b2(din_25_msk_ab2), .msk_a0b3(din_25_msk_ab3),
           .msk_a0b0_1sc(din_25_msk_ab0_1sc), .msk_a0b1_1sc(din_25_msk_ab1_1sc), .msk_a0b2_1sc(din_25_msk_ab2_1sc), .msk_a0b3_1sc(din_25_msk_ab3_1sc),

           .a1b0(din_27_ab0), .a1b1(din_27_ab1), .a1b2(din_27_ab2),
           .a1b0_1sc(din_27_ab0_1sc), .a1b1_1sc(din_27_ab1_1sc), .a1b2_1sc(din_27_ab2_1sc),
           .msk_a1b0(din_27_msk_ab0), .msk_a1b1(din_27_msk_ab1), .msk_a1b2(din_27_msk_ab2),
           .msk_a1b0_1sc(din_27_msk_ab0_1sc), .msk_a1b1_1sc(din_27_msk_ab1_1sc), .msk_a1b2_1sc(din_27_msk_ab2_1sc),

           .a2b0(din_29_ab0), .a2b1(din_29_ab1),
           .a2b0_1sc(din_29_ab0_1sc), .a2b1_1sc(din_29_ab1_1sc),
           .msk_a2b0(din_29_msk_ab0), .msk_a2b1(din_29_msk_ab1),
           .msk_a2b0_1sc(din_29_msk_ab0_1sc), .msk_a2b1_1sc(din_29_msk_ab1_1sc),
           
           .a3b0(din_31_ab0),
           .a3b0_1sc(din_31_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_26_calc (
           .clk(clk), .sign(din_signs_reg[26]), 
           .p(addr_0_26),
           .a0b0(din_26_ab0), .a0b1(din_26_ab1), .a0b2(din_26_ab2), .a0b3(din_26_ab3),
           .a0b0_1sc(din_26_ab0_1sc), .a0b1_1sc(din_26_ab1_1sc), .a0b2_1sc(din_26_ab2_1sc), .a0b3_1sc(din_26_ab3_1sc),
           .msk_a0b0(din_26_msk_ab0), .msk_a0b1(din_26_msk_ab1), .msk_a0b2(din_26_msk_ab2), .msk_a0b3(din_26_msk_ab3),
           .msk_a0b0_1sc(din_26_msk_ab0_1sc), .msk_a0b1_1sc(din_26_msk_ab1_1sc), .msk_a0b2_1sc(din_26_msk_ab2_1sc), .msk_a0b3_1sc(din_26_msk_ab3_1sc),

           .a1b0(din_28_ab0), .a1b1(din_28_ab1), .a1b2(din_28_ab2),
           .a1b0_1sc(din_28_ab0_1sc), .a1b1_1sc(din_28_ab1_1sc), .a1b2_1sc(din_28_ab2_1sc),
           .msk_a1b0(din_28_msk_ab0), .msk_a1b1(din_28_msk_ab1), .msk_a1b2(din_28_msk_ab2),
           .msk_a1b0_1sc(din_28_msk_ab0_1sc), .msk_a1b1_1sc(din_28_msk_ab1_1sc), .msk_a1b2_1sc(din_28_msk_ab2_1sc),

           .a2b0(din_30_ab0), .a2b1(din_30_ab1),
           .a2b0_1sc(din_30_ab0_1sc), .a2b1_1sc(din_30_ab1_1sc),
           .msk_a2b0(din_30_msk_ab0), .msk_a2b1(din_30_msk_ab1),
           .msk_a2b0_1sc(din_30_msk_ab0_1sc), .msk_a2b1_1sc(din_30_msk_ab1_1sc),
           
           .a3b0(din_32_ab0),
           .a3b0_1sc(din_32_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_27_calc (
           .clk(clk), .sign(din_signs_reg[27]), 
           .p(addr_0_27),
           .a0b0(din_27_ab0), .a0b1(din_27_ab1), .a0b2(din_27_ab2), .a0b3(din_27_ab3),
           .a0b0_1sc(din_27_ab0_1sc), .a0b1_1sc(din_27_ab1_1sc), .a0b2_1sc(din_27_ab2_1sc), .a0b3_1sc(din_27_ab3_1sc),
           .msk_a0b0(din_27_msk_ab0), .msk_a0b1(din_27_msk_ab1), .msk_a0b2(din_27_msk_ab2), .msk_a0b3(din_27_msk_ab3),
           .msk_a0b0_1sc(din_27_msk_ab0_1sc), .msk_a0b1_1sc(din_27_msk_ab1_1sc), .msk_a0b2_1sc(din_27_msk_ab2_1sc), .msk_a0b3_1sc(din_27_msk_ab3_1sc),

           .a1b0(din_29_ab0), .a1b1(din_29_ab1), .a1b2(din_29_ab2),
           .a1b0_1sc(din_29_ab0_1sc), .a1b1_1sc(din_29_ab1_1sc), .a1b2_1sc(din_29_ab2_1sc),
           .msk_a1b0(din_29_msk_ab0), .msk_a1b1(din_29_msk_ab1), .msk_a1b2(din_29_msk_ab2),
           .msk_a1b0_1sc(din_29_msk_ab0_1sc), .msk_a1b1_1sc(din_29_msk_ab1_1sc), .msk_a1b2_1sc(din_29_msk_ab2_1sc),

           .a2b0(din_31_ab0), .a2b1(din_31_ab1),
           .a2b0_1sc(din_31_ab0_1sc), .a2b1_1sc(din_31_ab1_1sc),
           .msk_a2b0(din_31_msk_ab0), .msk_a2b1(din_31_msk_ab1),
           .msk_a2b0_1sc(din_31_msk_ab0_1sc), .msk_a2b1_1sc(din_31_msk_ab1_1sc),
           
           .a3b0(din_33_ab0),
           .a3b0_1sc(din_33_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_28_calc (
           .clk(clk), .sign(din_signs_reg[28]), 
           .p(addr_0_28),
           .a0b0(din_28_ab0), .a0b1(din_28_ab1), .a0b2(din_28_ab2), .a0b3(din_28_ab3),
           .a0b0_1sc(din_28_ab0_1sc), .a0b1_1sc(din_28_ab1_1sc), .a0b2_1sc(din_28_ab2_1sc), .a0b3_1sc(din_28_ab3_1sc),
           .msk_a0b0(din_28_msk_ab0), .msk_a0b1(din_28_msk_ab1), .msk_a0b2(din_28_msk_ab2), .msk_a0b3(din_28_msk_ab3),
           .msk_a0b0_1sc(din_28_msk_ab0_1sc), .msk_a0b1_1sc(din_28_msk_ab1_1sc), .msk_a0b2_1sc(din_28_msk_ab2_1sc), .msk_a0b3_1sc(din_28_msk_ab3_1sc),

           .a1b0(din_30_ab0), .a1b1(din_30_ab1), .a1b2(din_30_ab2),
           .a1b0_1sc(din_30_ab0_1sc), .a1b1_1sc(din_30_ab1_1sc), .a1b2_1sc(din_30_ab2_1sc),
           .msk_a1b0(din_30_msk_ab0), .msk_a1b1(din_30_msk_ab1), .msk_a1b2(din_30_msk_ab2),
           .msk_a1b0_1sc(din_30_msk_ab0_1sc), .msk_a1b1_1sc(din_30_msk_ab1_1sc), .msk_a1b2_1sc(din_30_msk_ab2_1sc),

           .a2b0(din_32_ab0), .a2b1(din_32_ab1),
           .a2b0_1sc(din_32_ab0_1sc), .a2b1_1sc(din_32_ab1_1sc),
           .msk_a2b0(din_32_msk_ab0), .msk_a2b1(din_32_msk_ab1),
           .msk_a2b0_1sc(din_32_msk_ab0_1sc), .msk_a2b1_1sc(din_32_msk_ab1_1sc),
           
           .a3b0(din_34_ab0),
           .a3b0_1sc(din_34_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_29_calc (
           .clk(clk), .sign(din_signs_reg[29]), 
           .p(addr_0_29),
           .a0b0(din_29_ab0), .a0b1(din_29_ab1), .a0b2(din_29_ab2), .a0b3(din_29_ab3),
           .a0b0_1sc(din_29_ab0_1sc), .a0b1_1sc(din_29_ab1_1sc), .a0b2_1sc(din_29_ab2_1sc), .a0b3_1sc(din_29_ab3_1sc),
           .msk_a0b0(din_29_msk_ab0), .msk_a0b1(din_29_msk_ab1), .msk_a0b2(din_29_msk_ab2), .msk_a0b3(din_29_msk_ab3),
           .msk_a0b0_1sc(din_29_msk_ab0_1sc), .msk_a0b1_1sc(din_29_msk_ab1_1sc), .msk_a0b2_1sc(din_29_msk_ab2_1sc), .msk_a0b3_1sc(din_29_msk_ab3_1sc),

           .a1b0(din_31_ab0), .a1b1(din_31_ab1), .a1b2(din_31_ab2),
           .a1b0_1sc(din_31_ab0_1sc), .a1b1_1sc(din_31_ab1_1sc), .a1b2_1sc(din_31_ab2_1sc),
           .msk_a1b0(din_31_msk_ab0), .msk_a1b1(din_31_msk_ab1), .msk_a1b2(din_31_msk_ab2),
           .msk_a1b0_1sc(din_31_msk_ab0_1sc), .msk_a1b1_1sc(din_31_msk_ab1_1sc), .msk_a1b2_1sc(din_31_msk_ab2_1sc),

           .a2b0(din_33_ab0), .a2b1(din_33_ab1),
           .a2b0_1sc(din_33_ab0_1sc), .a2b1_1sc(din_33_ab1_1sc),
           .msk_a2b0(din_33_msk_ab0), .msk_a2b1(din_33_msk_ab1),
           .msk_a2b0_1sc(din_33_msk_ab0_1sc), .msk_a2b1_1sc(din_33_msk_ab1_1sc),
           
           .a3b0(din_35_ab0),
           .a3b0_1sc(din_35_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_30_calc (
           .clk(clk), .sign(din_signs_reg[30]), 
           .p(addr_0_30),
           .a0b0(din_30_ab0), .a0b1(din_30_ab1), .a0b2(din_30_ab2), .a0b3(din_30_ab3),
           .a0b0_1sc(din_30_ab0_1sc), .a0b1_1sc(din_30_ab1_1sc), .a0b2_1sc(din_30_ab2_1sc), .a0b3_1sc(din_30_ab3_1sc),
           .msk_a0b0(din_30_msk_ab0), .msk_a0b1(din_30_msk_ab1), .msk_a0b2(din_30_msk_ab2), .msk_a0b3(din_30_msk_ab3),
           .msk_a0b0_1sc(din_30_msk_ab0_1sc), .msk_a0b1_1sc(din_30_msk_ab1_1sc), .msk_a0b2_1sc(din_30_msk_ab2_1sc), .msk_a0b3_1sc(din_30_msk_ab3_1sc),

           .a1b0(din_32_ab0), .a1b1(din_32_ab1), .a1b2(din_32_ab2),
           .a1b0_1sc(din_32_ab0_1sc), .a1b1_1sc(din_32_ab1_1sc), .a1b2_1sc(din_32_ab2_1sc),
           .msk_a1b0(din_32_msk_ab0), .msk_a1b1(din_32_msk_ab1), .msk_a1b2(din_32_msk_ab2),
           .msk_a1b0_1sc(din_32_msk_ab0_1sc), .msk_a1b1_1sc(din_32_msk_ab1_1sc), .msk_a1b2_1sc(din_32_msk_ab2_1sc),

           .a2b0(din_34_ab0), .a2b1(din_34_ab1),
           .a2b0_1sc(din_34_ab0_1sc), .a2b1_1sc(din_34_ab1_1sc),
           .msk_a2b0(din_34_msk_ab0), .msk_a2b1(din_34_msk_ab1),
           .msk_a2b0_1sc(din_34_msk_ab0_1sc), .msk_a2b1_1sc(din_34_msk_ab1_1sc),
           
           .a3b0(din_36_ab0),
           .a3b0_1sc(din_36_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_0_31_calc (
           .clk(clk), .sign(din_signs_reg[31]), 
           .p(addr_0_31),
           .a0b0(din_31_ab0), .a0b1(din_31_ab1), .a0b2(din_31_ab2), .a0b3(din_31_ab3),
           .a0b0_1sc(din_31_ab0_1sc), .a0b1_1sc(din_31_ab1_1sc), .a0b2_1sc(din_31_ab2_1sc), .a0b3_1sc(din_31_ab3_1sc),
           .msk_a0b0(din_31_msk_ab0), .msk_a0b1(din_31_msk_ab1), .msk_a0b2(din_31_msk_ab2), .msk_a0b3(din_31_msk_ab3),
           .msk_a0b0_1sc(din_31_msk_ab0_1sc), .msk_a0b1_1sc(din_31_msk_ab1_1sc), .msk_a0b2_1sc(din_31_msk_ab2_1sc), .msk_a0b3_1sc(din_31_msk_ab3_1sc),

           .a1b0(din_33_ab0), .a1b1(din_33_ab1), .a1b2(din_33_ab2),
           .a1b0_1sc(din_33_ab0_1sc), .a1b1_1sc(din_33_ab1_1sc), .a1b2_1sc(din_33_ab2_1sc),
           .msk_a1b0(din_33_msk_ab0), .msk_a1b1(din_33_msk_ab1), .msk_a1b2(din_33_msk_ab2),
           .msk_a1b0_1sc(din_33_msk_ab0_1sc), .msk_a1b1_1sc(din_33_msk_ab1_1sc), .msk_a1b2_1sc(din_33_msk_ab2_1sc),

           .a2b0(din_35_ab0), .a2b1(din_35_ab1),
           .a2b0_1sc(din_35_ab0_1sc), .a2b1_1sc(din_35_ab1_1sc),
           .msk_a2b0(din_35_msk_ab0), .msk_a2b1(din_35_msk_ab1),
           .msk_a2b0_1sc(din_35_msk_ab0_1sc), .msk_a2b1_1sc(din_35_msk_ab1_1sc),
           
           .a3b0(din_37_ab0),
           .a3b0_1sc(din_37_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_0_calc (
           .clk(clk), .sign(din_signs_reg[0]), 
           .p(addr_1_0),
           .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
           .a0b0_1sc(din_0_ab0_1sc), .a0b1_1sc(din_0_ab1_1sc), .a0b2_1sc(din_0_ab2_1sc), .a0b3_1sc(din_0_ab3_1sc),
           .msk_a0b0(din_0_msk_ab0), .msk_a0b1(din_0_msk_ab1), .msk_a0b2(din_0_msk_ab2), .msk_a0b3(din_0_msk_ab3),
           .msk_a0b0_1sc(din_0_msk_ab0_1sc), .msk_a0b1_1sc(din_0_msk_ab1_1sc), .msk_a0b2_1sc(din_0_msk_ab2_1sc), .msk_a0b3_1sc(din_0_msk_ab3_1sc),

           .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2),
           .a1b0_1sc(din_2_ab0_1sc), .a1b1_1sc(din_2_ab1_1sc), .a1b2_1sc(din_2_ab2_1sc),
           .msk_a1b0(din_2_msk_ab0), .msk_a1b1(din_2_msk_ab1), .msk_a1b2(din_2_msk_ab2),
           .msk_a1b0_1sc(din_2_msk_ab0_1sc), .msk_a1b1_1sc(din_2_msk_ab1_1sc), .msk_a1b2_1sc(din_2_msk_ab2_1sc),

           .a2b0(din_4_ab0), .a2b1(din_4_ab1),
           .a2b0_1sc(din_4_ab0_1sc), .a2b1_1sc(din_4_ab1_1sc),
           .msk_a2b0(din_4_msk_ab0), .msk_a2b1(din_4_msk_ab1),
           .msk_a2b0_1sc(din_4_msk_ab0_1sc), .msk_a2b1_1sc(din_4_msk_ab1_1sc),
           
           .a3b0(din_6_ab0),
           .a3b0_1sc(din_6_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_1_calc (
           .clk(clk), .sign(din_signs_reg[1]), 
           .p(addr_1_1),
           .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
           .a0b0_1sc(din_1_ab0_1sc), .a0b1_1sc(din_1_ab1_1sc), .a0b2_1sc(din_1_ab2_1sc), .a0b3_1sc(din_1_ab3_1sc),
           .msk_a0b0(din_1_msk_ab0), .msk_a0b1(din_1_msk_ab1), .msk_a0b2(din_1_msk_ab2), .msk_a0b3(din_1_msk_ab3),
           .msk_a0b0_1sc(din_1_msk_ab0_1sc), .msk_a0b1_1sc(din_1_msk_ab1_1sc), .msk_a0b2_1sc(din_1_msk_ab2_1sc), .msk_a0b3_1sc(din_1_msk_ab3_1sc),

           .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2),
           .a1b0_1sc(din_3_ab0_1sc), .a1b1_1sc(din_3_ab1_1sc), .a1b2_1sc(din_3_ab2_1sc),
           .msk_a1b0(din_3_msk_ab0), .msk_a1b1(din_3_msk_ab1), .msk_a1b2(din_3_msk_ab2),
           .msk_a1b0_1sc(din_3_msk_ab0_1sc), .msk_a1b1_1sc(din_3_msk_ab1_1sc), .msk_a1b2_1sc(din_3_msk_ab2_1sc),

           .a2b0(din_5_ab0), .a2b1(din_5_ab1),
           .a2b0_1sc(din_5_ab0_1sc), .a2b1_1sc(din_5_ab1_1sc),
           .msk_a2b0(din_5_msk_ab0), .msk_a2b1(din_5_msk_ab1),
           .msk_a2b0_1sc(din_5_msk_ab0_1sc), .msk_a2b1_1sc(din_5_msk_ab1_1sc),
           
           .a3b0(din_7_ab0),
           .a3b0_1sc(din_7_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_2_calc (
           .clk(clk), .sign(din_signs_reg[2]), 
           .p(addr_1_2),
           .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
           .a0b0_1sc(din_2_ab0_1sc), .a0b1_1sc(din_2_ab1_1sc), .a0b2_1sc(din_2_ab2_1sc), .a0b3_1sc(din_2_ab3_1sc),
           .msk_a0b0(din_2_msk_ab0), .msk_a0b1(din_2_msk_ab1), .msk_a0b2(din_2_msk_ab2), .msk_a0b3(din_2_msk_ab3),
           .msk_a0b0_1sc(din_2_msk_ab0_1sc), .msk_a0b1_1sc(din_2_msk_ab1_1sc), .msk_a0b2_1sc(din_2_msk_ab2_1sc), .msk_a0b3_1sc(din_2_msk_ab3_1sc),

           .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2),
           .a1b0_1sc(din_4_ab0_1sc), .a1b1_1sc(din_4_ab1_1sc), .a1b2_1sc(din_4_ab2_1sc),
           .msk_a1b0(din_4_msk_ab0), .msk_a1b1(din_4_msk_ab1), .msk_a1b2(din_4_msk_ab2),
           .msk_a1b0_1sc(din_4_msk_ab0_1sc), .msk_a1b1_1sc(din_4_msk_ab1_1sc), .msk_a1b2_1sc(din_4_msk_ab2_1sc),

           .a2b0(din_6_ab0), .a2b1(din_6_ab1),
           .a2b0_1sc(din_6_ab0_1sc), .a2b1_1sc(din_6_ab1_1sc),
           .msk_a2b0(din_6_msk_ab0), .msk_a2b1(din_6_msk_ab1),
           .msk_a2b0_1sc(din_6_msk_ab0_1sc), .msk_a2b1_1sc(din_6_msk_ab1_1sc),
           
           .a3b0(din_8_ab0),
           .a3b0_1sc(din_8_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_3_calc (
           .clk(clk), .sign(din_signs_reg[3]), 
           .p(addr_1_3),
           .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
           .a0b0_1sc(din_3_ab0_1sc), .a0b1_1sc(din_3_ab1_1sc), .a0b2_1sc(din_3_ab2_1sc), .a0b3_1sc(din_3_ab3_1sc),
           .msk_a0b0(din_3_msk_ab0), .msk_a0b1(din_3_msk_ab1), .msk_a0b2(din_3_msk_ab2), .msk_a0b3(din_3_msk_ab3),
           .msk_a0b0_1sc(din_3_msk_ab0_1sc), .msk_a0b1_1sc(din_3_msk_ab1_1sc), .msk_a0b2_1sc(din_3_msk_ab2_1sc), .msk_a0b3_1sc(din_3_msk_ab3_1sc),

           .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2),
           .a1b0_1sc(din_5_ab0_1sc), .a1b1_1sc(din_5_ab1_1sc), .a1b2_1sc(din_5_ab2_1sc),
           .msk_a1b0(din_5_msk_ab0), .msk_a1b1(din_5_msk_ab1), .msk_a1b2(din_5_msk_ab2),
           .msk_a1b0_1sc(din_5_msk_ab0_1sc), .msk_a1b1_1sc(din_5_msk_ab1_1sc), .msk_a1b2_1sc(din_5_msk_ab2_1sc),

           .a2b0(din_7_ab0), .a2b1(din_7_ab1),
           .a2b0_1sc(din_7_ab0_1sc), .a2b1_1sc(din_7_ab1_1sc),
           .msk_a2b0(din_7_msk_ab0), .msk_a2b1(din_7_msk_ab1),
           .msk_a2b0_1sc(din_7_msk_ab0_1sc), .msk_a2b1_1sc(din_7_msk_ab1_1sc),
           
           .a3b0(din_9_ab0),
           .a3b0_1sc(din_9_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_4_calc (
           .clk(clk), .sign(din_signs_reg[4]), 
           .p(addr_1_4),
           .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
           .a0b0_1sc(din_4_ab0_1sc), .a0b1_1sc(din_4_ab1_1sc), .a0b2_1sc(din_4_ab2_1sc), .a0b3_1sc(din_4_ab3_1sc),
           .msk_a0b0(din_4_msk_ab0), .msk_a0b1(din_4_msk_ab1), .msk_a0b2(din_4_msk_ab2), .msk_a0b3(din_4_msk_ab3),
           .msk_a0b0_1sc(din_4_msk_ab0_1sc), .msk_a0b1_1sc(din_4_msk_ab1_1sc), .msk_a0b2_1sc(din_4_msk_ab2_1sc), .msk_a0b3_1sc(din_4_msk_ab3_1sc),

           .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2),
           .a1b0_1sc(din_6_ab0_1sc), .a1b1_1sc(din_6_ab1_1sc), .a1b2_1sc(din_6_ab2_1sc),
           .msk_a1b0(din_6_msk_ab0), .msk_a1b1(din_6_msk_ab1), .msk_a1b2(din_6_msk_ab2),
           .msk_a1b0_1sc(din_6_msk_ab0_1sc), .msk_a1b1_1sc(din_6_msk_ab1_1sc), .msk_a1b2_1sc(din_6_msk_ab2_1sc),

           .a2b0(din_8_ab0), .a2b1(din_8_ab1),
           .a2b0_1sc(din_8_ab0_1sc), .a2b1_1sc(din_8_ab1_1sc),
           .msk_a2b0(din_8_msk_ab0), .msk_a2b1(din_8_msk_ab1),
           .msk_a2b0_1sc(din_8_msk_ab0_1sc), .msk_a2b1_1sc(din_8_msk_ab1_1sc),
           
           .a3b0(din_10_ab0),
           .a3b0_1sc(din_10_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_5_calc (
           .clk(clk), .sign(din_signs_reg[5]), 
           .p(addr_1_5),
           .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
           .a0b0_1sc(din_5_ab0_1sc), .a0b1_1sc(din_5_ab1_1sc), .a0b2_1sc(din_5_ab2_1sc), .a0b3_1sc(din_5_ab3_1sc),
           .msk_a0b0(din_5_msk_ab0), .msk_a0b1(din_5_msk_ab1), .msk_a0b2(din_5_msk_ab2), .msk_a0b3(din_5_msk_ab3),
           .msk_a0b0_1sc(din_5_msk_ab0_1sc), .msk_a0b1_1sc(din_5_msk_ab1_1sc), .msk_a0b2_1sc(din_5_msk_ab2_1sc), .msk_a0b3_1sc(din_5_msk_ab3_1sc),

           .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2),
           .a1b0_1sc(din_7_ab0_1sc), .a1b1_1sc(din_7_ab1_1sc), .a1b2_1sc(din_7_ab2_1sc),
           .msk_a1b0(din_7_msk_ab0), .msk_a1b1(din_7_msk_ab1), .msk_a1b2(din_7_msk_ab2),
           .msk_a1b0_1sc(din_7_msk_ab0_1sc), .msk_a1b1_1sc(din_7_msk_ab1_1sc), .msk_a1b2_1sc(din_7_msk_ab2_1sc),

           .a2b0(din_9_ab0), .a2b1(din_9_ab1),
           .a2b0_1sc(din_9_ab0_1sc), .a2b1_1sc(din_9_ab1_1sc),
           .msk_a2b0(din_9_msk_ab0), .msk_a2b1(din_9_msk_ab1),
           .msk_a2b0_1sc(din_9_msk_ab0_1sc), .msk_a2b1_1sc(din_9_msk_ab1_1sc),
           
           .a3b0(din_11_ab0),
           .a3b0_1sc(din_11_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_6_calc (
           .clk(clk), .sign(din_signs_reg[6]), 
           .p(addr_1_6),
           .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
           .a0b0_1sc(din_6_ab0_1sc), .a0b1_1sc(din_6_ab1_1sc), .a0b2_1sc(din_6_ab2_1sc), .a0b3_1sc(din_6_ab3_1sc),
           .msk_a0b0(din_6_msk_ab0), .msk_a0b1(din_6_msk_ab1), .msk_a0b2(din_6_msk_ab2), .msk_a0b3(din_6_msk_ab3),
           .msk_a0b0_1sc(din_6_msk_ab0_1sc), .msk_a0b1_1sc(din_6_msk_ab1_1sc), .msk_a0b2_1sc(din_6_msk_ab2_1sc), .msk_a0b3_1sc(din_6_msk_ab3_1sc),

           .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2),
           .a1b0_1sc(din_8_ab0_1sc), .a1b1_1sc(din_8_ab1_1sc), .a1b2_1sc(din_8_ab2_1sc),
           .msk_a1b0(din_8_msk_ab0), .msk_a1b1(din_8_msk_ab1), .msk_a1b2(din_8_msk_ab2),
           .msk_a1b0_1sc(din_8_msk_ab0_1sc), .msk_a1b1_1sc(din_8_msk_ab1_1sc), .msk_a1b2_1sc(din_8_msk_ab2_1sc),

           .a2b0(din_10_ab0), .a2b1(din_10_ab1),
           .a2b0_1sc(din_10_ab0_1sc), .a2b1_1sc(din_10_ab1_1sc),
           .msk_a2b0(din_10_msk_ab0), .msk_a2b1(din_10_msk_ab1),
           .msk_a2b0_1sc(din_10_msk_ab0_1sc), .msk_a2b1_1sc(din_10_msk_ab1_1sc),
           
           .a3b0(din_12_ab0),
           .a3b0_1sc(din_12_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_7_calc (
           .clk(clk), .sign(din_signs_reg[7]), 
           .p(addr_1_7),
           .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
           .a0b0_1sc(din_7_ab0_1sc), .a0b1_1sc(din_7_ab1_1sc), .a0b2_1sc(din_7_ab2_1sc), .a0b3_1sc(din_7_ab3_1sc),
           .msk_a0b0(din_7_msk_ab0), .msk_a0b1(din_7_msk_ab1), .msk_a0b2(din_7_msk_ab2), .msk_a0b3(din_7_msk_ab3),
           .msk_a0b0_1sc(din_7_msk_ab0_1sc), .msk_a0b1_1sc(din_7_msk_ab1_1sc), .msk_a0b2_1sc(din_7_msk_ab2_1sc), .msk_a0b3_1sc(din_7_msk_ab3_1sc),

           .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2),
           .a1b0_1sc(din_9_ab0_1sc), .a1b1_1sc(din_9_ab1_1sc), .a1b2_1sc(din_9_ab2_1sc),
           .msk_a1b0(din_9_msk_ab0), .msk_a1b1(din_9_msk_ab1), .msk_a1b2(din_9_msk_ab2),
           .msk_a1b0_1sc(din_9_msk_ab0_1sc), .msk_a1b1_1sc(din_9_msk_ab1_1sc), .msk_a1b2_1sc(din_9_msk_ab2_1sc),

           .a2b0(din_11_ab0), .a2b1(din_11_ab1),
           .a2b0_1sc(din_11_ab0_1sc), .a2b1_1sc(din_11_ab1_1sc),
           .msk_a2b0(din_11_msk_ab0), .msk_a2b1(din_11_msk_ab1),
           .msk_a2b0_1sc(din_11_msk_ab0_1sc), .msk_a2b1_1sc(din_11_msk_ab1_1sc),
           
           .a3b0(din_13_ab0),
           .a3b0_1sc(din_13_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_8_calc (
           .clk(clk), .sign(din_signs_reg[8]), 
           .p(addr_1_8),
           .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
           .a0b0_1sc(din_8_ab0_1sc), .a0b1_1sc(din_8_ab1_1sc), .a0b2_1sc(din_8_ab2_1sc), .a0b3_1sc(din_8_ab3_1sc),
           .msk_a0b0(din_8_msk_ab0), .msk_a0b1(din_8_msk_ab1), .msk_a0b2(din_8_msk_ab2), .msk_a0b3(din_8_msk_ab3),
           .msk_a0b0_1sc(din_8_msk_ab0_1sc), .msk_a0b1_1sc(din_8_msk_ab1_1sc), .msk_a0b2_1sc(din_8_msk_ab2_1sc), .msk_a0b3_1sc(din_8_msk_ab3_1sc),

           .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2),
           .a1b0_1sc(din_10_ab0_1sc), .a1b1_1sc(din_10_ab1_1sc), .a1b2_1sc(din_10_ab2_1sc),
           .msk_a1b0(din_10_msk_ab0), .msk_a1b1(din_10_msk_ab1), .msk_a1b2(din_10_msk_ab2),
           .msk_a1b0_1sc(din_10_msk_ab0_1sc), .msk_a1b1_1sc(din_10_msk_ab1_1sc), .msk_a1b2_1sc(din_10_msk_ab2_1sc),

           .a2b0(din_12_ab0), .a2b1(din_12_ab1),
           .a2b0_1sc(din_12_ab0_1sc), .a2b1_1sc(din_12_ab1_1sc),
           .msk_a2b0(din_12_msk_ab0), .msk_a2b1(din_12_msk_ab1),
           .msk_a2b0_1sc(din_12_msk_ab0_1sc), .msk_a2b1_1sc(din_12_msk_ab1_1sc),
           
           .a3b0(din_14_ab0),
           .a3b0_1sc(din_14_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_9_calc (
           .clk(clk), .sign(din_signs_reg[9]), 
           .p(addr_1_9),
           .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
           .a0b0_1sc(din_9_ab0_1sc), .a0b1_1sc(din_9_ab1_1sc), .a0b2_1sc(din_9_ab2_1sc), .a0b3_1sc(din_9_ab3_1sc),
           .msk_a0b0(din_9_msk_ab0), .msk_a0b1(din_9_msk_ab1), .msk_a0b2(din_9_msk_ab2), .msk_a0b3(din_9_msk_ab3),
           .msk_a0b0_1sc(din_9_msk_ab0_1sc), .msk_a0b1_1sc(din_9_msk_ab1_1sc), .msk_a0b2_1sc(din_9_msk_ab2_1sc), .msk_a0b3_1sc(din_9_msk_ab3_1sc),

           .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2),
           .a1b0_1sc(din_11_ab0_1sc), .a1b1_1sc(din_11_ab1_1sc), .a1b2_1sc(din_11_ab2_1sc),
           .msk_a1b0(din_11_msk_ab0), .msk_a1b1(din_11_msk_ab1), .msk_a1b2(din_11_msk_ab2),
           .msk_a1b0_1sc(din_11_msk_ab0_1sc), .msk_a1b1_1sc(din_11_msk_ab1_1sc), .msk_a1b2_1sc(din_11_msk_ab2_1sc),

           .a2b0(din_13_ab0), .a2b1(din_13_ab1),
           .a2b0_1sc(din_13_ab0_1sc), .a2b1_1sc(din_13_ab1_1sc),
           .msk_a2b0(din_13_msk_ab0), .msk_a2b1(din_13_msk_ab1),
           .msk_a2b0_1sc(din_13_msk_ab0_1sc), .msk_a2b1_1sc(din_13_msk_ab1_1sc),
           
           .a3b0(din_15_ab0),
           .a3b0_1sc(din_15_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_10_calc (
           .clk(clk), .sign(din_signs_reg[10]), 
           .p(addr_1_10),
           .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
           .a0b0_1sc(din_10_ab0_1sc), .a0b1_1sc(din_10_ab1_1sc), .a0b2_1sc(din_10_ab2_1sc), .a0b3_1sc(din_10_ab3_1sc),
           .msk_a0b0(din_10_msk_ab0), .msk_a0b1(din_10_msk_ab1), .msk_a0b2(din_10_msk_ab2), .msk_a0b3(din_10_msk_ab3),
           .msk_a0b0_1sc(din_10_msk_ab0_1sc), .msk_a0b1_1sc(din_10_msk_ab1_1sc), .msk_a0b2_1sc(din_10_msk_ab2_1sc), .msk_a0b3_1sc(din_10_msk_ab3_1sc),

           .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2),
           .a1b0_1sc(din_12_ab0_1sc), .a1b1_1sc(din_12_ab1_1sc), .a1b2_1sc(din_12_ab2_1sc),
           .msk_a1b0(din_12_msk_ab0), .msk_a1b1(din_12_msk_ab1), .msk_a1b2(din_12_msk_ab2),
           .msk_a1b0_1sc(din_12_msk_ab0_1sc), .msk_a1b1_1sc(din_12_msk_ab1_1sc), .msk_a1b2_1sc(din_12_msk_ab2_1sc),

           .a2b0(din_14_ab0), .a2b1(din_14_ab1),
           .a2b0_1sc(din_14_ab0_1sc), .a2b1_1sc(din_14_ab1_1sc),
           .msk_a2b0(din_14_msk_ab0), .msk_a2b1(din_14_msk_ab1),
           .msk_a2b0_1sc(din_14_msk_ab0_1sc), .msk_a2b1_1sc(din_14_msk_ab1_1sc),
           
           .a3b0(din_16_ab0),
           .a3b0_1sc(din_16_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_11_calc (
           .clk(clk), .sign(din_signs_reg[11]), 
           .p(addr_1_11),
           .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
           .a0b0_1sc(din_11_ab0_1sc), .a0b1_1sc(din_11_ab1_1sc), .a0b2_1sc(din_11_ab2_1sc), .a0b3_1sc(din_11_ab3_1sc),
           .msk_a0b0(din_11_msk_ab0), .msk_a0b1(din_11_msk_ab1), .msk_a0b2(din_11_msk_ab2), .msk_a0b3(din_11_msk_ab3),
           .msk_a0b0_1sc(din_11_msk_ab0_1sc), .msk_a0b1_1sc(din_11_msk_ab1_1sc), .msk_a0b2_1sc(din_11_msk_ab2_1sc), .msk_a0b3_1sc(din_11_msk_ab3_1sc),

           .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2),
           .a1b0_1sc(din_13_ab0_1sc), .a1b1_1sc(din_13_ab1_1sc), .a1b2_1sc(din_13_ab2_1sc),
           .msk_a1b0(din_13_msk_ab0), .msk_a1b1(din_13_msk_ab1), .msk_a1b2(din_13_msk_ab2),
           .msk_a1b0_1sc(din_13_msk_ab0_1sc), .msk_a1b1_1sc(din_13_msk_ab1_1sc), .msk_a1b2_1sc(din_13_msk_ab2_1sc),

           .a2b0(din_15_ab0), .a2b1(din_15_ab1),
           .a2b0_1sc(din_15_ab0_1sc), .a2b1_1sc(din_15_ab1_1sc),
           .msk_a2b0(din_15_msk_ab0), .msk_a2b1(din_15_msk_ab1),
           .msk_a2b0_1sc(din_15_msk_ab0_1sc), .msk_a2b1_1sc(din_15_msk_ab1_1sc),
           
           .a3b0(din_17_ab0),
           .a3b0_1sc(din_17_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_12_calc (
           .clk(clk), .sign(din_signs_reg[12]), 
           .p(addr_1_12),
           .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
           .a0b0_1sc(din_12_ab0_1sc), .a0b1_1sc(din_12_ab1_1sc), .a0b2_1sc(din_12_ab2_1sc), .a0b3_1sc(din_12_ab3_1sc),
           .msk_a0b0(din_12_msk_ab0), .msk_a0b1(din_12_msk_ab1), .msk_a0b2(din_12_msk_ab2), .msk_a0b3(din_12_msk_ab3),
           .msk_a0b0_1sc(din_12_msk_ab0_1sc), .msk_a0b1_1sc(din_12_msk_ab1_1sc), .msk_a0b2_1sc(din_12_msk_ab2_1sc), .msk_a0b3_1sc(din_12_msk_ab3_1sc),

           .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2),
           .a1b0_1sc(din_14_ab0_1sc), .a1b1_1sc(din_14_ab1_1sc), .a1b2_1sc(din_14_ab2_1sc),
           .msk_a1b0(din_14_msk_ab0), .msk_a1b1(din_14_msk_ab1), .msk_a1b2(din_14_msk_ab2),
           .msk_a1b0_1sc(din_14_msk_ab0_1sc), .msk_a1b1_1sc(din_14_msk_ab1_1sc), .msk_a1b2_1sc(din_14_msk_ab2_1sc),

           .a2b0(din_16_ab0), .a2b1(din_16_ab1),
           .a2b0_1sc(din_16_ab0_1sc), .a2b1_1sc(din_16_ab1_1sc),
           .msk_a2b0(din_16_msk_ab0), .msk_a2b1(din_16_msk_ab1),
           .msk_a2b0_1sc(din_16_msk_ab0_1sc), .msk_a2b1_1sc(din_16_msk_ab1_1sc),
           
           .a3b0(din_18_ab0),
           .a3b0_1sc(din_18_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_13_calc (
           .clk(clk), .sign(din_signs_reg[13]), 
           .p(addr_1_13),
           .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
           .a0b0_1sc(din_13_ab0_1sc), .a0b1_1sc(din_13_ab1_1sc), .a0b2_1sc(din_13_ab2_1sc), .a0b3_1sc(din_13_ab3_1sc),
           .msk_a0b0(din_13_msk_ab0), .msk_a0b1(din_13_msk_ab1), .msk_a0b2(din_13_msk_ab2), .msk_a0b3(din_13_msk_ab3),
           .msk_a0b0_1sc(din_13_msk_ab0_1sc), .msk_a0b1_1sc(din_13_msk_ab1_1sc), .msk_a0b2_1sc(din_13_msk_ab2_1sc), .msk_a0b3_1sc(din_13_msk_ab3_1sc),

           .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2),
           .a1b0_1sc(din_15_ab0_1sc), .a1b1_1sc(din_15_ab1_1sc), .a1b2_1sc(din_15_ab2_1sc),
           .msk_a1b0(din_15_msk_ab0), .msk_a1b1(din_15_msk_ab1), .msk_a1b2(din_15_msk_ab2),
           .msk_a1b0_1sc(din_15_msk_ab0_1sc), .msk_a1b1_1sc(din_15_msk_ab1_1sc), .msk_a1b2_1sc(din_15_msk_ab2_1sc),

           .a2b0(din_17_ab0), .a2b1(din_17_ab1),
           .a2b0_1sc(din_17_ab0_1sc), .a2b1_1sc(din_17_ab1_1sc),
           .msk_a2b0(din_17_msk_ab0), .msk_a2b1(din_17_msk_ab1),
           .msk_a2b0_1sc(din_17_msk_ab0_1sc), .msk_a2b1_1sc(din_17_msk_ab1_1sc),
           
           .a3b0(din_19_ab0),
           .a3b0_1sc(din_19_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_14_calc (
           .clk(clk), .sign(din_signs_reg[14]), 
           .p(addr_1_14),
           .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
           .a0b0_1sc(din_14_ab0_1sc), .a0b1_1sc(din_14_ab1_1sc), .a0b2_1sc(din_14_ab2_1sc), .a0b3_1sc(din_14_ab3_1sc),
           .msk_a0b0(din_14_msk_ab0), .msk_a0b1(din_14_msk_ab1), .msk_a0b2(din_14_msk_ab2), .msk_a0b3(din_14_msk_ab3),
           .msk_a0b0_1sc(din_14_msk_ab0_1sc), .msk_a0b1_1sc(din_14_msk_ab1_1sc), .msk_a0b2_1sc(din_14_msk_ab2_1sc), .msk_a0b3_1sc(din_14_msk_ab3_1sc),

           .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2),
           .a1b0_1sc(din_16_ab0_1sc), .a1b1_1sc(din_16_ab1_1sc), .a1b2_1sc(din_16_ab2_1sc),
           .msk_a1b0(din_16_msk_ab0), .msk_a1b1(din_16_msk_ab1), .msk_a1b2(din_16_msk_ab2),
           .msk_a1b0_1sc(din_16_msk_ab0_1sc), .msk_a1b1_1sc(din_16_msk_ab1_1sc), .msk_a1b2_1sc(din_16_msk_ab2_1sc),

           .a2b0(din_18_ab0), .a2b1(din_18_ab1),
           .a2b0_1sc(din_18_ab0_1sc), .a2b1_1sc(din_18_ab1_1sc),
           .msk_a2b0(din_18_msk_ab0), .msk_a2b1(din_18_msk_ab1),
           .msk_a2b0_1sc(din_18_msk_ab0_1sc), .msk_a2b1_1sc(din_18_msk_ab1_1sc),
           
           .a3b0(din_20_ab0),
           .a3b0_1sc(din_20_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_15_calc (
           .clk(clk), .sign(din_signs_reg[15]), 
           .p(addr_1_15),
           .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
           .a0b0_1sc(din_15_ab0_1sc), .a0b1_1sc(din_15_ab1_1sc), .a0b2_1sc(din_15_ab2_1sc), .a0b3_1sc(din_15_ab3_1sc),
           .msk_a0b0(din_15_msk_ab0), .msk_a0b1(din_15_msk_ab1), .msk_a0b2(din_15_msk_ab2), .msk_a0b3(din_15_msk_ab3),
           .msk_a0b0_1sc(din_15_msk_ab0_1sc), .msk_a0b1_1sc(din_15_msk_ab1_1sc), .msk_a0b2_1sc(din_15_msk_ab2_1sc), .msk_a0b3_1sc(din_15_msk_ab3_1sc),

           .a1b0(din_17_ab0), .a1b1(din_17_ab1), .a1b2(din_17_ab2),
           .a1b0_1sc(din_17_ab0_1sc), .a1b1_1sc(din_17_ab1_1sc), .a1b2_1sc(din_17_ab2_1sc),
           .msk_a1b0(din_17_msk_ab0), .msk_a1b1(din_17_msk_ab1), .msk_a1b2(din_17_msk_ab2),
           .msk_a1b0_1sc(din_17_msk_ab0_1sc), .msk_a1b1_1sc(din_17_msk_ab1_1sc), .msk_a1b2_1sc(din_17_msk_ab2_1sc),

           .a2b0(din_19_ab0), .a2b1(din_19_ab1),
           .a2b0_1sc(din_19_ab0_1sc), .a2b1_1sc(din_19_ab1_1sc),
           .msk_a2b0(din_19_msk_ab0), .msk_a2b1(din_19_msk_ab1),
           .msk_a2b0_1sc(din_19_msk_ab0_1sc), .msk_a2b1_1sc(din_19_msk_ab1_1sc),
           
           .a3b0(din_21_ab0),
           .a3b0_1sc(din_21_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_16_calc (
           .clk(clk), .sign(din_signs_reg[16]), 
           .p(addr_1_16),
           .a0b0(din_16_ab0), .a0b1(din_16_ab1), .a0b2(din_16_ab2), .a0b3(din_16_ab3),
           .a0b0_1sc(din_16_ab0_1sc), .a0b1_1sc(din_16_ab1_1sc), .a0b2_1sc(din_16_ab2_1sc), .a0b3_1sc(din_16_ab3_1sc),
           .msk_a0b0(din_16_msk_ab0), .msk_a0b1(din_16_msk_ab1), .msk_a0b2(din_16_msk_ab2), .msk_a0b3(din_16_msk_ab3),
           .msk_a0b0_1sc(din_16_msk_ab0_1sc), .msk_a0b1_1sc(din_16_msk_ab1_1sc), .msk_a0b2_1sc(din_16_msk_ab2_1sc), .msk_a0b3_1sc(din_16_msk_ab3_1sc),

           .a1b0(din_18_ab0), .a1b1(din_18_ab1), .a1b2(din_18_ab2),
           .a1b0_1sc(din_18_ab0_1sc), .a1b1_1sc(din_18_ab1_1sc), .a1b2_1sc(din_18_ab2_1sc),
           .msk_a1b0(din_18_msk_ab0), .msk_a1b1(din_18_msk_ab1), .msk_a1b2(din_18_msk_ab2),
           .msk_a1b0_1sc(din_18_msk_ab0_1sc), .msk_a1b1_1sc(din_18_msk_ab1_1sc), .msk_a1b2_1sc(din_18_msk_ab2_1sc),

           .a2b0(din_20_ab0), .a2b1(din_20_ab1),
           .a2b0_1sc(din_20_ab0_1sc), .a2b1_1sc(din_20_ab1_1sc),
           .msk_a2b0(din_20_msk_ab0), .msk_a2b1(din_20_msk_ab1),
           .msk_a2b0_1sc(din_20_msk_ab0_1sc), .msk_a2b1_1sc(din_20_msk_ab1_1sc),
           
           .a3b0(din_22_ab0),
           .a3b0_1sc(din_22_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_17_calc (
           .clk(clk), .sign(din_signs_reg[17]), 
           .p(addr_1_17),
           .a0b0(din_17_ab0), .a0b1(din_17_ab1), .a0b2(din_17_ab2), .a0b3(din_17_ab3),
           .a0b0_1sc(din_17_ab0_1sc), .a0b1_1sc(din_17_ab1_1sc), .a0b2_1sc(din_17_ab2_1sc), .a0b3_1sc(din_17_ab3_1sc),
           .msk_a0b0(din_17_msk_ab0), .msk_a0b1(din_17_msk_ab1), .msk_a0b2(din_17_msk_ab2), .msk_a0b3(din_17_msk_ab3),
           .msk_a0b0_1sc(din_17_msk_ab0_1sc), .msk_a0b1_1sc(din_17_msk_ab1_1sc), .msk_a0b2_1sc(din_17_msk_ab2_1sc), .msk_a0b3_1sc(din_17_msk_ab3_1sc),

           .a1b0(din_19_ab0), .a1b1(din_19_ab1), .a1b2(din_19_ab2),
           .a1b0_1sc(din_19_ab0_1sc), .a1b1_1sc(din_19_ab1_1sc), .a1b2_1sc(din_19_ab2_1sc),
           .msk_a1b0(din_19_msk_ab0), .msk_a1b1(din_19_msk_ab1), .msk_a1b2(din_19_msk_ab2),
           .msk_a1b0_1sc(din_19_msk_ab0_1sc), .msk_a1b1_1sc(din_19_msk_ab1_1sc), .msk_a1b2_1sc(din_19_msk_ab2_1sc),

           .a2b0(din_21_ab0), .a2b1(din_21_ab1),
           .a2b0_1sc(din_21_ab0_1sc), .a2b1_1sc(din_21_ab1_1sc),
           .msk_a2b0(din_21_msk_ab0), .msk_a2b1(din_21_msk_ab1),
           .msk_a2b0_1sc(din_21_msk_ab0_1sc), .msk_a2b1_1sc(din_21_msk_ab1_1sc),
           
           .a3b0(din_23_ab0),
           .a3b0_1sc(din_23_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_18_calc (
           .clk(clk), .sign(din_signs_reg[18]), 
           .p(addr_1_18),
           .a0b0(din_18_ab0), .a0b1(din_18_ab1), .a0b2(din_18_ab2), .a0b3(din_18_ab3),
           .a0b0_1sc(din_18_ab0_1sc), .a0b1_1sc(din_18_ab1_1sc), .a0b2_1sc(din_18_ab2_1sc), .a0b3_1sc(din_18_ab3_1sc),
           .msk_a0b0(din_18_msk_ab0), .msk_a0b1(din_18_msk_ab1), .msk_a0b2(din_18_msk_ab2), .msk_a0b3(din_18_msk_ab3),
           .msk_a0b0_1sc(din_18_msk_ab0_1sc), .msk_a0b1_1sc(din_18_msk_ab1_1sc), .msk_a0b2_1sc(din_18_msk_ab2_1sc), .msk_a0b3_1sc(din_18_msk_ab3_1sc),

           .a1b0(din_20_ab0), .a1b1(din_20_ab1), .a1b2(din_20_ab2),
           .a1b0_1sc(din_20_ab0_1sc), .a1b1_1sc(din_20_ab1_1sc), .a1b2_1sc(din_20_ab2_1sc),
           .msk_a1b0(din_20_msk_ab0), .msk_a1b1(din_20_msk_ab1), .msk_a1b2(din_20_msk_ab2),
           .msk_a1b0_1sc(din_20_msk_ab0_1sc), .msk_a1b1_1sc(din_20_msk_ab1_1sc), .msk_a1b2_1sc(din_20_msk_ab2_1sc),

           .a2b0(din_22_ab0), .a2b1(din_22_ab1),
           .a2b0_1sc(din_22_ab0_1sc), .a2b1_1sc(din_22_ab1_1sc),
           .msk_a2b0(din_22_msk_ab0), .msk_a2b1(din_22_msk_ab1),
           .msk_a2b0_1sc(din_22_msk_ab0_1sc), .msk_a2b1_1sc(din_22_msk_ab1_1sc),
           
           .a3b0(din_24_ab0),
           .a3b0_1sc(din_24_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_19_calc (
           .clk(clk), .sign(din_signs_reg[19]), 
           .p(addr_1_19),
           .a0b0(din_19_ab0), .a0b1(din_19_ab1), .a0b2(din_19_ab2), .a0b3(din_19_ab3),
           .a0b0_1sc(din_19_ab0_1sc), .a0b1_1sc(din_19_ab1_1sc), .a0b2_1sc(din_19_ab2_1sc), .a0b3_1sc(din_19_ab3_1sc),
           .msk_a0b0(din_19_msk_ab0), .msk_a0b1(din_19_msk_ab1), .msk_a0b2(din_19_msk_ab2), .msk_a0b3(din_19_msk_ab3),
           .msk_a0b0_1sc(din_19_msk_ab0_1sc), .msk_a0b1_1sc(din_19_msk_ab1_1sc), .msk_a0b2_1sc(din_19_msk_ab2_1sc), .msk_a0b3_1sc(din_19_msk_ab3_1sc),

           .a1b0(din_21_ab0), .a1b1(din_21_ab1), .a1b2(din_21_ab2),
           .a1b0_1sc(din_21_ab0_1sc), .a1b1_1sc(din_21_ab1_1sc), .a1b2_1sc(din_21_ab2_1sc),
           .msk_a1b0(din_21_msk_ab0), .msk_a1b1(din_21_msk_ab1), .msk_a1b2(din_21_msk_ab2),
           .msk_a1b0_1sc(din_21_msk_ab0_1sc), .msk_a1b1_1sc(din_21_msk_ab1_1sc), .msk_a1b2_1sc(din_21_msk_ab2_1sc),

           .a2b0(din_23_ab0), .a2b1(din_23_ab1),
           .a2b0_1sc(din_23_ab0_1sc), .a2b1_1sc(din_23_ab1_1sc),
           .msk_a2b0(din_23_msk_ab0), .msk_a2b1(din_23_msk_ab1),
           .msk_a2b0_1sc(din_23_msk_ab0_1sc), .msk_a2b1_1sc(din_23_msk_ab1_1sc),
           
           .a3b0(din_25_ab0),
           .a3b0_1sc(din_25_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_20_calc (
           .clk(clk), .sign(din_signs_reg[20]), 
           .p(addr_1_20),
           .a0b0(din_20_ab0), .a0b1(din_20_ab1), .a0b2(din_20_ab2), .a0b3(din_20_ab3),
           .a0b0_1sc(din_20_ab0_1sc), .a0b1_1sc(din_20_ab1_1sc), .a0b2_1sc(din_20_ab2_1sc), .a0b3_1sc(din_20_ab3_1sc),
           .msk_a0b0(din_20_msk_ab0), .msk_a0b1(din_20_msk_ab1), .msk_a0b2(din_20_msk_ab2), .msk_a0b3(din_20_msk_ab3),
           .msk_a0b0_1sc(din_20_msk_ab0_1sc), .msk_a0b1_1sc(din_20_msk_ab1_1sc), .msk_a0b2_1sc(din_20_msk_ab2_1sc), .msk_a0b3_1sc(din_20_msk_ab3_1sc),

           .a1b0(din_22_ab0), .a1b1(din_22_ab1), .a1b2(din_22_ab2),
           .a1b0_1sc(din_22_ab0_1sc), .a1b1_1sc(din_22_ab1_1sc), .a1b2_1sc(din_22_ab2_1sc),
           .msk_a1b0(din_22_msk_ab0), .msk_a1b1(din_22_msk_ab1), .msk_a1b2(din_22_msk_ab2),
           .msk_a1b0_1sc(din_22_msk_ab0_1sc), .msk_a1b1_1sc(din_22_msk_ab1_1sc), .msk_a1b2_1sc(din_22_msk_ab2_1sc),

           .a2b0(din_24_ab0), .a2b1(din_24_ab1),
           .a2b0_1sc(din_24_ab0_1sc), .a2b1_1sc(din_24_ab1_1sc),
           .msk_a2b0(din_24_msk_ab0), .msk_a2b1(din_24_msk_ab1),
           .msk_a2b0_1sc(din_24_msk_ab0_1sc), .msk_a2b1_1sc(din_24_msk_ab1_1sc),
           
           .a3b0(din_26_ab0),
           .a3b0_1sc(din_26_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_21_calc (
           .clk(clk), .sign(din_signs_reg[21]), 
           .p(addr_1_21),
           .a0b0(din_21_ab0), .a0b1(din_21_ab1), .a0b2(din_21_ab2), .a0b3(din_21_ab3),
           .a0b0_1sc(din_21_ab0_1sc), .a0b1_1sc(din_21_ab1_1sc), .a0b2_1sc(din_21_ab2_1sc), .a0b3_1sc(din_21_ab3_1sc),
           .msk_a0b0(din_21_msk_ab0), .msk_a0b1(din_21_msk_ab1), .msk_a0b2(din_21_msk_ab2), .msk_a0b3(din_21_msk_ab3),
           .msk_a0b0_1sc(din_21_msk_ab0_1sc), .msk_a0b1_1sc(din_21_msk_ab1_1sc), .msk_a0b2_1sc(din_21_msk_ab2_1sc), .msk_a0b3_1sc(din_21_msk_ab3_1sc),

           .a1b0(din_23_ab0), .a1b1(din_23_ab1), .a1b2(din_23_ab2),
           .a1b0_1sc(din_23_ab0_1sc), .a1b1_1sc(din_23_ab1_1sc), .a1b2_1sc(din_23_ab2_1sc),
           .msk_a1b0(din_23_msk_ab0), .msk_a1b1(din_23_msk_ab1), .msk_a1b2(din_23_msk_ab2),
           .msk_a1b0_1sc(din_23_msk_ab0_1sc), .msk_a1b1_1sc(din_23_msk_ab1_1sc), .msk_a1b2_1sc(din_23_msk_ab2_1sc),

           .a2b0(din_25_ab0), .a2b1(din_25_ab1),
           .a2b0_1sc(din_25_ab0_1sc), .a2b1_1sc(din_25_ab1_1sc),
           .msk_a2b0(din_25_msk_ab0), .msk_a2b1(din_25_msk_ab1),
           .msk_a2b0_1sc(din_25_msk_ab0_1sc), .msk_a2b1_1sc(din_25_msk_ab1_1sc),
           
           .a3b0(din_27_ab0),
           .a3b0_1sc(din_27_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_22_calc (
           .clk(clk), .sign(din_signs_reg[22]), 
           .p(addr_1_22),
           .a0b0(din_22_ab0), .a0b1(din_22_ab1), .a0b2(din_22_ab2), .a0b3(din_22_ab3),
           .a0b0_1sc(din_22_ab0_1sc), .a0b1_1sc(din_22_ab1_1sc), .a0b2_1sc(din_22_ab2_1sc), .a0b3_1sc(din_22_ab3_1sc),
           .msk_a0b0(din_22_msk_ab0), .msk_a0b1(din_22_msk_ab1), .msk_a0b2(din_22_msk_ab2), .msk_a0b3(din_22_msk_ab3),
           .msk_a0b0_1sc(din_22_msk_ab0_1sc), .msk_a0b1_1sc(din_22_msk_ab1_1sc), .msk_a0b2_1sc(din_22_msk_ab2_1sc), .msk_a0b3_1sc(din_22_msk_ab3_1sc),

           .a1b0(din_24_ab0), .a1b1(din_24_ab1), .a1b2(din_24_ab2),
           .a1b0_1sc(din_24_ab0_1sc), .a1b1_1sc(din_24_ab1_1sc), .a1b2_1sc(din_24_ab2_1sc),
           .msk_a1b0(din_24_msk_ab0), .msk_a1b1(din_24_msk_ab1), .msk_a1b2(din_24_msk_ab2),
           .msk_a1b0_1sc(din_24_msk_ab0_1sc), .msk_a1b1_1sc(din_24_msk_ab1_1sc), .msk_a1b2_1sc(din_24_msk_ab2_1sc),

           .a2b0(din_26_ab0), .a2b1(din_26_ab1),
           .a2b0_1sc(din_26_ab0_1sc), .a2b1_1sc(din_26_ab1_1sc),
           .msk_a2b0(din_26_msk_ab0), .msk_a2b1(din_26_msk_ab1),
           .msk_a2b0_1sc(din_26_msk_ab0_1sc), .msk_a2b1_1sc(din_26_msk_ab1_1sc),
           
           .a3b0(din_28_ab0),
           .a3b0_1sc(din_28_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_23_calc (
           .clk(clk), .sign(din_signs_reg[23]), 
           .p(addr_1_23),
           .a0b0(din_23_ab0), .a0b1(din_23_ab1), .a0b2(din_23_ab2), .a0b3(din_23_ab3),
           .a0b0_1sc(din_23_ab0_1sc), .a0b1_1sc(din_23_ab1_1sc), .a0b2_1sc(din_23_ab2_1sc), .a0b3_1sc(din_23_ab3_1sc),
           .msk_a0b0(din_23_msk_ab0), .msk_a0b1(din_23_msk_ab1), .msk_a0b2(din_23_msk_ab2), .msk_a0b3(din_23_msk_ab3),
           .msk_a0b0_1sc(din_23_msk_ab0_1sc), .msk_a0b1_1sc(din_23_msk_ab1_1sc), .msk_a0b2_1sc(din_23_msk_ab2_1sc), .msk_a0b3_1sc(din_23_msk_ab3_1sc),

           .a1b0(din_25_ab0), .a1b1(din_25_ab1), .a1b2(din_25_ab2),
           .a1b0_1sc(din_25_ab0_1sc), .a1b1_1sc(din_25_ab1_1sc), .a1b2_1sc(din_25_ab2_1sc),
           .msk_a1b0(din_25_msk_ab0), .msk_a1b1(din_25_msk_ab1), .msk_a1b2(din_25_msk_ab2),
           .msk_a1b0_1sc(din_25_msk_ab0_1sc), .msk_a1b1_1sc(din_25_msk_ab1_1sc), .msk_a1b2_1sc(din_25_msk_ab2_1sc),

           .a2b0(din_27_ab0), .a2b1(din_27_ab1),
           .a2b0_1sc(din_27_ab0_1sc), .a2b1_1sc(din_27_ab1_1sc),
           .msk_a2b0(din_27_msk_ab0), .msk_a2b1(din_27_msk_ab1),
           .msk_a2b0_1sc(din_27_msk_ab0_1sc), .msk_a2b1_1sc(din_27_msk_ab1_1sc),
           
           .a3b0(din_29_ab0),
           .a3b0_1sc(din_29_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_24_calc (
           .clk(clk), .sign(din_signs_reg[24]), 
           .p(addr_1_24),
           .a0b0(din_24_ab0), .a0b1(din_24_ab1), .a0b2(din_24_ab2), .a0b3(din_24_ab3),
           .a0b0_1sc(din_24_ab0_1sc), .a0b1_1sc(din_24_ab1_1sc), .a0b2_1sc(din_24_ab2_1sc), .a0b3_1sc(din_24_ab3_1sc),
           .msk_a0b0(din_24_msk_ab0), .msk_a0b1(din_24_msk_ab1), .msk_a0b2(din_24_msk_ab2), .msk_a0b3(din_24_msk_ab3),
           .msk_a0b0_1sc(din_24_msk_ab0_1sc), .msk_a0b1_1sc(din_24_msk_ab1_1sc), .msk_a0b2_1sc(din_24_msk_ab2_1sc), .msk_a0b3_1sc(din_24_msk_ab3_1sc),

           .a1b0(din_26_ab0), .a1b1(din_26_ab1), .a1b2(din_26_ab2),
           .a1b0_1sc(din_26_ab0_1sc), .a1b1_1sc(din_26_ab1_1sc), .a1b2_1sc(din_26_ab2_1sc),
           .msk_a1b0(din_26_msk_ab0), .msk_a1b1(din_26_msk_ab1), .msk_a1b2(din_26_msk_ab2),
           .msk_a1b0_1sc(din_26_msk_ab0_1sc), .msk_a1b1_1sc(din_26_msk_ab1_1sc), .msk_a1b2_1sc(din_26_msk_ab2_1sc),

           .a2b0(din_28_ab0), .a2b1(din_28_ab1),
           .a2b0_1sc(din_28_ab0_1sc), .a2b1_1sc(din_28_ab1_1sc),
           .msk_a2b0(din_28_msk_ab0), .msk_a2b1(din_28_msk_ab1),
           .msk_a2b0_1sc(din_28_msk_ab0_1sc), .msk_a2b1_1sc(din_28_msk_ab1_1sc),
           
           .a3b0(din_30_ab0),
           .a3b0_1sc(din_30_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_25_calc (
           .clk(clk), .sign(din_signs_reg[25]), 
           .p(addr_1_25),
           .a0b0(din_25_ab0), .a0b1(din_25_ab1), .a0b2(din_25_ab2), .a0b3(din_25_ab3),
           .a0b0_1sc(din_25_ab0_1sc), .a0b1_1sc(din_25_ab1_1sc), .a0b2_1sc(din_25_ab2_1sc), .a0b3_1sc(din_25_ab3_1sc),
           .msk_a0b0(din_25_msk_ab0), .msk_a0b1(din_25_msk_ab1), .msk_a0b2(din_25_msk_ab2), .msk_a0b3(din_25_msk_ab3),
           .msk_a0b0_1sc(din_25_msk_ab0_1sc), .msk_a0b1_1sc(din_25_msk_ab1_1sc), .msk_a0b2_1sc(din_25_msk_ab2_1sc), .msk_a0b3_1sc(din_25_msk_ab3_1sc),

           .a1b0(din_27_ab0), .a1b1(din_27_ab1), .a1b2(din_27_ab2),
           .a1b0_1sc(din_27_ab0_1sc), .a1b1_1sc(din_27_ab1_1sc), .a1b2_1sc(din_27_ab2_1sc),
           .msk_a1b0(din_27_msk_ab0), .msk_a1b1(din_27_msk_ab1), .msk_a1b2(din_27_msk_ab2),
           .msk_a1b0_1sc(din_27_msk_ab0_1sc), .msk_a1b1_1sc(din_27_msk_ab1_1sc), .msk_a1b2_1sc(din_27_msk_ab2_1sc),

           .a2b0(din_29_ab0), .a2b1(din_29_ab1),
           .a2b0_1sc(din_29_ab0_1sc), .a2b1_1sc(din_29_ab1_1sc),
           .msk_a2b0(din_29_msk_ab0), .msk_a2b1(din_29_msk_ab1),
           .msk_a2b0_1sc(din_29_msk_ab0_1sc), .msk_a2b1_1sc(din_29_msk_ab1_1sc),
           
           .a3b0(din_31_ab0),
           .a3b0_1sc(din_31_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_26_calc (
           .clk(clk), .sign(din_signs_reg[26]), 
           .p(addr_1_26),
           .a0b0(din_26_ab0), .a0b1(din_26_ab1), .a0b2(din_26_ab2), .a0b3(din_26_ab3),
           .a0b0_1sc(din_26_ab0_1sc), .a0b1_1sc(din_26_ab1_1sc), .a0b2_1sc(din_26_ab2_1sc), .a0b3_1sc(din_26_ab3_1sc),
           .msk_a0b0(din_26_msk_ab0), .msk_a0b1(din_26_msk_ab1), .msk_a0b2(din_26_msk_ab2), .msk_a0b3(din_26_msk_ab3),
           .msk_a0b0_1sc(din_26_msk_ab0_1sc), .msk_a0b1_1sc(din_26_msk_ab1_1sc), .msk_a0b2_1sc(din_26_msk_ab2_1sc), .msk_a0b3_1sc(din_26_msk_ab3_1sc),

           .a1b0(din_28_ab0), .a1b1(din_28_ab1), .a1b2(din_28_ab2),
           .a1b0_1sc(din_28_ab0_1sc), .a1b1_1sc(din_28_ab1_1sc), .a1b2_1sc(din_28_ab2_1sc),
           .msk_a1b0(din_28_msk_ab0), .msk_a1b1(din_28_msk_ab1), .msk_a1b2(din_28_msk_ab2),
           .msk_a1b0_1sc(din_28_msk_ab0_1sc), .msk_a1b1_1sc(din_28_msk_ab1_1sc), .msk_a1b2_1sc(din_28_msk_ab2_1sc),

           .a2b0(din_30_ab0), .a2b1(din_30_ab1),
           .a2b0_1sc(din_30_ab0_1sc), .a2b1_1sc(din_30_ab1_1sc),
           .msk_a2b0(din_30_msk_ab0), .msk_a2b1(din_30_msk_ab1),
           .msk_a2b0_1sc(din_30_msk_ab0_1sc), .msk_a2b1_1sc(din_30_msk_ab1_1sc),
           
           .a3b0(din_32_ab0),
           .a3b0_1sc(din_32_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_27_calc (
           .clk(clk), .sign(din_signs_reg[27]), 
           .p(addr_1_27),
           .a0b0(din_27_ab0), .a0b1(din_27_ab1), .a0b2(din_27_ab2), .a0b3(din_27_ab3),
           .a0b0_1sc(din_27_ab0_1sc), .a0b1_1sc(din_27_ab1_1sc), .a0b2_1sc(din_27_ab2_1sc), .a0b3_1sc(din_27_ab3_1sc),
           .msk_a0b0(din_27_msk_ab0), .msk_a0b1(din_27_msk_ab1), .msk_a0b2(din_27_msk_ab2), .msk_a0b3(din_27_msk_ab3),
           .msk_a0b0_1sc(din_27_msk_ab0_1sc), .msk_a0b1_1sc(din_27_msk_ab1_1sc), .msk_a0b2_1sc(din_27_msk_ab2_1sc), .msk_a0b3_1sc(din_27_msk_ab3_1sc),

           .a1b0(din_29_ab0), .a1b1(din_29_ab1), .a1b2(din_29_ab2),
           .a1b0_1sc(din_29_ab0_1sc), .a1b1_1sc(din_29_ab1_1sc), .a1b2_1sc(din_29_ab2_1sc),
           .msk_a1b0(din_29_msk_ab0), .msk_a1b1(din_29_msk_ab1), .msk_a1b2(din_29_msk_ab2),
           .msk_a1b0_1sc(din_29_msk_ab0_1sc), .msk_a1b1_1sc(din_29_msk_ab1_1sc), .msk_a1b2_1sc(din_29_msk_ab2_1sc),

           .a2b0(din_31_ab0), .a2b1(din_31_ab1),
           .a2b0_1sc(din_31_ab0_1sc), .a2b1_1sc(din_31_ab1_1sc),
           .msk_a2b0(din_31_msk_ab0), .msk_a2b1(din_31_msk_ab1),
           .msk_a2b0_1sc(din_31_msk_ab0_1sc), .msk_a2b1_1sc(din_31_msk_ab1_1sc),
           
           .a3b0(din_33_ab0),
           .a3b0_1sc(din_33_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_28_calc (
           .clk(clk), .sign(din_signs_reg[28]), 
           .p(addr_1_28),
           .a0b0(din_28_ab0), .a0b1(din_28_ab1), .a0b2(din_28_ab2), .a0b3(din_28_ab3),
           .a0b0_1sc(din_28_ab0_1sc), .a0b1_1sc(din_28_ab1_1sc), .a0b2_1sc(din_28_ab2_1sc), .a0b3_1sc(din_28_ab3_1sc),
           .msk_a0b0(din_28_msk_ab0), .msk_a0b1(din_28_msk_ab1), .msk_a0b2(din_28_msk_ab2), .msk_a0b3(din_28_msk_ab3),
           .msk_a0b0_1sc(din_28_msk_ab0_1sc), .msk_a0b1_1sc(din_28_msk_ab1_1sc), .msk_a0b2_1sc(din_28_msk_ab2_1sc), .msk_a0b3_1sc(din_28_msk_ab3_1sc),

           .a1b0(din_30_ab0), .a1b1(din_30_ab1), .a1b2(din_30_ab2),
           .a1b0_1sc(din_30_ab0_1sc), .a1b1_1sc(din_30_ab1_1sc), .a1b2_1sc(din_30_ab2_1sc),
           .msk_a1b0(din_30_msk_ab0), .msk_a1b1(din_30_msk_ab1), .msk_a1b2(din_30_msk_ab2),
           .msk_a1b0_1sc(din_30_msk_ab0_1sc), .msk_a1b1_1sc(din_30_msk_ab1_1sc), .msk_a1b2_1sc(din_30_msk_ab2_1sc),

           .a2b0(din_32_ab0), .a2b1(din_32_ab1),
           .a2b0_1sc(din_32_ab0_1sc), .a2b1_1sc(din_32_ab1_1sc),
           .msk_a2b0(din_32_msk_ab0), .msk_a2b1(din_32_msk_ab1),
           .msk_a2b0_1sc(din_32_msk_ab0_1sc), .msk_a2b1_1sc(din_32_msk_ab1_1sc),
           
           .a3b0(din_34_ab0),
           .a3b0_1sc(din_34_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_29_calc (
           .clk(clk), .sign(din_signs_reg[29]), 
           .p(addr_1_29),
           .a0b0(din_29_ab0), .a0b1(din_29_ab1), .a0b2(din_29_ab2), .a0b3(din_29_ab3),
           .a0b0_1sc(din_29_ab0_1sc), .a0b1_1sc(din_29_ab1_1sc), .a0b2_1sc(din_29_ab2_1sc), .a0b3_1sc(din_29_ab3_1sc),
           .msk_a0b0(din_29_msk_ab0), .msk_a0b1(din_29_msk_ab1), .msk_a0b2(din_29_msk_ab2), .msk_a0b3(din_29_msk_ab3),
           .msk_a0b0_1sc(din_29_msk_ab0_1sc), .msk_a0b1_1sc(din_29_msk_ab1_1sc), .msk_a0b2_1sc(din_29_msk_ab2_1sc), .msk_a0b3_1sc(din_29_msk_ab3_1sc),

           .a1b0(din_31_ab0), .a1b1(din_31_ab1), .a1b2(din_31_ab2),
           .a1b0_1sc(din_31_ab0_1sc), .a1b1_1sc(din_31_ab1_1sc), .a1b2_1sc(din_31_ab2_1sc),
           .msk_a1b0(din_31_msk_ab0), .msk_a1b1(din_31_msk_ab1), .msk_a1b2(din_31_msk_ab2),
           .msk_a1b0_1sc(din_31_msk_ab0_1sc), .msk_a1b1_1sc(din_31_msk_ab1_1sc), .msk_a1b2_1sc(din_31_msk_ab2_1sc),

           .a2b0(din_33_ab0), .a2b1(din_33_ab1),
           .a2b0_1sc(din_33_ab0_1sc), .a2b1_1sc(din_33_ab1_1sc),
           .msk_a2b0(din_33_msk_ab0), .msk_a2b1(din_33_msk_ab1),
           .msk_a2b0_1sc(din_33_msk_ab0_1sc), .msk_a2b1_1sc(din_33_msk_ab1_1sc),
           
           .a3b0(din_35_ab0),
           .a3b0_1sc(din_35_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_30_calc (
           .clk(clk), .sign(din_signs_reg[30]), 
           .p(addr_1_30),
           .a0b0(din_30_ab0), .a0b1(din_30_ab1), .a0b2(din_30_ab2), .a0b3(din_30_ab3),
           .a0b0_1sc(din_30_ab0_1sc), .a0b1_1sc(din_30_ab1_1sc), .a0b2_1sc(din_30_ab2_1sc), .a0b3_1sc(din_30_ab3_1sc),
           .msk_a0b0(din_30_msk_ab0), .msk_a0b1(din_30_msk_ab1), .msk_a0b2(din_30_msk_ab2), .msk_a0b3(din_30_msk_ab3),
           .msk_a0b0_1sc(din_30_msk_ab0_1sc), .msk_a0b1_1sc(din_30_msk_ab1_1sc), .msk_a0b2_1sc(din_30_msk_ab2_1sc), .msk_a0b3_1sc(din_30_msk_ab3_1sc),

           .a1b0(din_32_ab0), .a1b1(din_32_ab1), .a1b2(din_32_ab2),
           .a1b0_1sc(din_32_ab0_1sc), .a1b1_1sc(din_32_ab1_1sc), .a1b2_1sc(din_32_ab2_1sc),
           .msk_a1b0(din_32_msk_ab0), .msk_a1b1(din_32_msk_ab1), .msk_a1b2(din_32_msk_ab2),
           .msk_a1b0_1sc(din_32_msk_ab0_1sc), .msk_a1b1_1sc(din_32_msk_ab1_1sc), .msk_a1b2_1sc(din_32_msk_ab2_1sc),

           .a2b0(din_34_ab0), .a2b1(din_34_ab1),
           .a2b0_1sc(din_34_ab0_1sc), .a2b1_1sc(din_34_ab1_1sc),
           .msk_a2b0(din_34_msk_ab0), .msk_a2b1(din_34_msk_ab1),
           .msk_a2b0_1sc(din_34_msk_ab0_1sc), .msk_a2b1_1sc(din_34_msk_ab1_1sc),
           
           .a3b0(din_36_ab0),
           .a3b0_1sc(din_36_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15)
) addr_1_31_calc (
           .clk(clk), .sign(din_signs_reg[31]), 
           .p(addr_1_31),
           .a0b0(din_31_ab0), .a0b1(din_31_ab1), .a0b2(din_31_ab2), .a0b3(din_31_ab3),
           .a0b0_1sc(din_31_ab0_1sc), .a0b1_1sc(din_31_ab1_1sc), .a0b2_1sc(din_31_ab2_1sc), .a0b3_1sc(din_31_ab3_1sc),
           .msk_a0b0(din_31_msk_ab0), .msk_a0b1(din_31_msk_ab1), .msk_a0b2(din_31_msk_ab2), .msk_a0b3(din_31_msk_ab3),
           .msk_a0b0_1sc(din_31_msk_ab0_1sc), .msk_a0b1_1sc(din_31_msk_ab1_1sc), .msk_a0b2_1sc(din_31_msk_ab2_1sc), .msk_a0b3_1sc(din_31_msk_ab3_1sc),

           .a1b0(din_33_ab0), .a1b1(din_33_ab1), .a1b2(din_33_ab2),
           .a1b0_1sc(din_33_ab0_1sc), .a1b1_1sc(din_33_ab1_1sc), .a1b2_1sc(din_33_ab2_1sc),
           .msk_a1b0(din_33_msk_ab0), .msk_a1b1(din_33_msk_ab1), .msk_a1b2(din_33_msk_ab2),
           .msk_a1b0_1sc(din_33_msk_ab0_1sc), .msk_a1b1_1sc(din_33_msk_ab1_1sc), .msk_a1b2_1sc(din_33_msk_ab2_1sc),

           .a2b0(din_35_ab0), .a2b1(din_35_ab1),
           .a2b0_1sc(din_35_ab0_1sc), .a2b1_1sc(din_35_ab1_1sc),
           .msk_a2b0(din_35_msk_ab0), .msk_a2b1(din_35_msk_ab1),
           .msk_a2b0_1sc(din_35_msk_ab0_1sc), .msk_a2b1_1sc(din_35_msk_ab1_1sc),
           
           .a3b0(din_37_ab0),
           .a3b0_1sc(din_37_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_0_calc (
           .clk(clk), .sign(din_signs_reg[0]), 
           .p(addr_2_0),
           .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
           .a0b0_1sc(din_0_ab0_1sc), .a0b1_1sc(din_0_ab1_1sc), .a0b2_1sc(din_0_ab2_1sc), .a0b3_1sc(din_0_ab3_1sc),
           .msk_a0b0(din_0_msk_ab0), .msk_a0b1(din_0_msk_ab1), .msk_a0b2(din_0_msk_ab2), .msk_a0b3(din_0_msk_ab3),
           .msk_a0b0_1sc(din_0_msk_ab0_1sc), .msk_a0b1_1sc(din_0_msk_ab1_1sc), .msk_a0b2_1sc(din_0_msk_ab2_1sc), .msk_a0b3_1sc(din_0_msk_ab3_1sc),

           .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2),
           .a1b0_1sc(din_2_ab0_1sc), .a1b1_1sc(din_2_ab1_1sc), .a1b2_1sc(din_2_ab2_1sc),
           .msk_a1b0(din_2_msk_ab0), .msk_a1b1(din_2_msk_ab1), .msk_a1b2(din_2_msk_ab2),
           .msk_a1b0_1sc(din_2_msk_ab0_1sc), .msk_a1b1_1sc(din_2_msk_ab1_1sc), .msk_a1b2_1sc(din_2_msk_ab2_1sc),

           .a2b0(din_4_ab0), .a2b1(din_4_ab1),
           .a2b0_1sc(din_4_ab0_1sc), .a2b1_1sc(din_4_ab1_1sc),
           .msk_a2b0(din_4_msk_ab0), .msk_a2b1(din_4_msk_ab1),
           .msk_a2b0_1sc(din_4_msk_ab0_1sc), .msk_a2b1_1sc(din_4_msk_ab1_1sc),
           
           .a3b0(din_6_ab0),
           .a3b0_1sc(din_6_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_1_calc (
           .clk(clk), .sign(din_signs_reg[1]), 
           .p(addr_2_1),
           .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
           .a0b0_1sc(din_1_ab0_1sc), .a0b1_1sc(din_1_ab1_1sc), .a0b2_1sc(din_1_ab2_1sc), .a0b3_1sc(din_1_ab3_1sc),
           .msk_a0b0(din_1_msk_ab0), .msk_a0b1(din_1_msk_ab1), .msk_a0b2(din_1_msk_ab2), .msk_a0b3(din_1_msk_ab3),
           .msk_a0b0_1sc(din_1_msk_ab0_1sc), .msk_a0b1_1sc(din_1_msk_ab1_1sc), .msk_a0b2_1sc(din_1_msk_ab2_1sc), .msk_a0b3_1sc(din_1_msk_ab3_1sc),

           .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2),
           .a1b0_1sc(din_3_ab0_1sc), .a1b1_1sc(din_3_ab1_1sc), .a1b2_1sc(din_3_ab2_1sc),
           .msk_a1b0(din_3_msk_ab0), .msk_a1b1(din_3_msk_ab1), .msk_a1b2(din_3_msk_ab2),
           .msk_a1b0_1sc(din_3_msk_ab0_1sc), .msk_a1b1_1sc(din_3_msk_ab1_1sc), .msk_a1b2_1sc(din_3_msk_ab2_1sc),

           .a2b0(din_5_ab0), .a2b1(din_5_ab1),
           .a2b0_1sc(din_5_ab0_1sc), .a2b1_1sc(din_5_ab1_1sc),
           .msk_a2b0(din_5_msk_ab0), .msk_a2b1(din_5_msk_ab1),
           .msk_a2b0_1sc(din_5_msk_ab0_1sc), .msk_a2b1_1sc(din_5_msk_ab1_1sc),
           
           .a3b0(din_7_ab0),
           .a3b0_1sc(din_7_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_2_calc (
           .clk(clk), .sign(din_signs_reg[2]), 
           .p(addr_2_2),
           .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
           .a0b0_1sc(din_2_ab0_1sc), .a0b1_1sc(din_2_ab1_1sc), .a0b2_1sc(din_2_ab2_1sc), .a0b3_1sc(din_2_ab3_1sc),
           .msk_a0b0(din_2_msk_ab0), .msk_a0b1(din_2_msk_ab1), .msk_a0b2(din_2_msk_ab2), .msk_a0b3(din_2_msk_ab3),
           .msk_a0b0_1sc(din_2_msk_ab0_1sc), .msk_a0b1_1sc(din_2_msk_ab1_1sc), .msk_a0b2_1sc(din_2_msk_ab2_1sc), .msk_a0b3_1sc(din_2_msk_ab3_1sc),

           .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2),
           .a1b0_1sc(din_4_ab0_1sc), .a1b1_1sc(din_4_ab1_1sc), .a1b2_1sc(din_4_ab2_1sc),
           .msk_a1b0(din_4_msk_ab0), .msk_a1b1(din_4_msk_ab1), .msk_a1b2(din_4_msk_ab2),
           .msk_a1b0_1sc(din_4_msk_ab0_1sc), .msk_a1b1_1sc(din_4_msk_ab1_1sc), .msk_a1b2_1sc(din_4_msk_ab2_1sc),

           .a2b0(din_6_ab0), .a2b1(din_6_ab1),
           .a2b0_1sc(din_6_ab0_1sc), .a2b1_1sc(din_6_ab1_1sc),
           .msk_a2b0(din_6_msk_ab0), .msk_a2b1(din_6_msk_ab1),
           .msk_a2b0_1sc(din_6_msk_ab0_1sc), .msk_a2b1_1sc(din_6_msk_ab1_1sc),
           
           .a3b0(din_8_ab0),
           .a3b0_1sc(din_8_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_3_calc (
           .clk(clk), .sign(din_signs_reg[3]), 
           .p(addr_2_3),
           .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
           .a0b0_1sc(din_3_ab0_1sc), .a0b1_1sc(din_3_ab1_1sc), .a0b2_1sc(din_3_ab2_1sc), .a0b3_1sc(din_3_ab3_1sc),
           .msk_a0b0(din_3_msk_ab0), .msk_a0b1(din_3_msk_ab1), .msk_a0b2(din_3_msk_ab2), .msk_a0b3(din_3_msk_ab3),
           .msk_a0b0_1sc(din_3_msk_ab0_1sc), .msk_a0b1_1sc(din_3_msk_ab1_1sc), .msk_a0b2_1sc(din_3_msk_ab2_1sc), .msk_a0b3_1sc(din_3_msk_ab3_1sc),

           .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2),
           .a1b0_1sc(din_5_ab0_1sc), .a1b1_1sc(din_5_ab1_1sc), .a1b2_1sc(din_5_ab2_1sc),
           .msk_a1b0(din_5_msk_ab0), .msk_a1b1(din_5_msk_ab1), .msk_a1b2(din_5_msk_ab2),
           .msk_a1b0_1sc(din_5_msk_ab0_1sc), .msk_a1b1_1sc(din_5_msk_ab1_1sc), .msk_a1b2_1sc(din_5_msk_ab2_1sc),

           .a2b0(din_7_ab0), .a2b1(din_7_ab1),
           .a2b0_1sc(din_7_ab0_1sc), .a2b1_1sc(din_7_ab1_1sc),
           .msk_a2b0(din_7_msk_ab0), .msk_a2b1(din_7_msk_ab1),
           .msk_a2b0_1sc(din_7_msk_ab0_1sc), .msk_a2b1_1sc(din_7_msk_ab1_1sc),
           
           .a3b0(din_9_ab0),
           .a3b0_1sc(din_9_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_4_calc (
           .clk(clk), .sign(din_signs_reg[4]), 
           .p(addr_2_4),
           .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
           .a0b0_1sc(din_4_ab0_1sc), .a0b1_1sc(din_4_ab1_1sc), .a0b2_1sc(din_4_ab2_1sc), .a0b3_1sc(din_4_ab3_1sc),
           .msk_a0b0(din_4_msk_ab0), .msk_a0b1(din_4_msk_ab1), .msk_a0b2(din_4_msk_ab2), .msk_a0b3(din_4_msk_ab3),
           .msk_a0b0_1sc(din_4_msk_ab0_1sc), .msk_a0b1_1sc(din_4_msk_ab1_1sc), .msk_a0b2_1sc(din_4_msk_ab2_1sc), .msk_a0b3_1sc(din_4_msk_ab3_1sc),

           .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2),
           .a1b0_1sc(din_6_ab0_1sc), .a1b1_1sc(din_6_ab1_1sc), .a1b2_1sc(din_6_ab2_1sc),
           .msk_a1b0(din_6_msk_ab0), .msk_a1b1(din_6_msk_ab1), .msk_a1b2(din_6_msk_ab2),
           .msk_a1b0_1sc(din_6_msk_ab0_1sc), .msk_a1b1_1sc(din_6_msk_ab1_1sc), .msk_a1b2_1sc(din_6_msk_ab2_1sc),

           .a2b0(din_8_ab0), .a2b1(din_8_ab1),
           .a2b0_1sc(din_8_ab0_1sc), .a2b1_1sc(din_8_ab1_1sc),
           .msk_a2b0(din_8_msk_ab0), .msk_a2b1(din_8_msk_ab1),
           .msk_a2b0_1sc(din_8_msk_ab0_1sc), .msk_a2b1_1sc(din_8_msk_ab1_1sc),
           
           .a3b0(din_10_ab0),
           .a3b0_1sc(din_10_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_5_calc (
           .clk(clk), .sign(din_signs_reg[5]), 
           .p(addr_2_5),
           .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
           .a0b0_1sc(din_5_ab0_1sc), .a0b1_1sc(din_5_ab1_1sc), .a0b2_1sc(din_5_ab2_1sc), .a0b3_1sc(din_5_ab3_1sc),
           .msk_a0b0(din_5_msk_ab0), .msk_a0b1(din_5_msk_ab1), .msk_a0b2(din_5_msk_ab2), .msk_a0b3(din_5_msk_ab3),
           .msk_a0b0_1sc(din_5_msk_ab0_1sc), .msk_a0b1_1sc(din_5_msk_ab1_1sc), .msk_a0b2_1sc(din_5_msk_ab2_1sc), .msk_a0b3_1sc(din_5_msk_ab3_1sc),

           .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2),
           .a1b0_1sc(din_7_ab0_1sc), .a1b1_1sc(din_7_ab1_1sc), .a1b2_1sc(din_7_ab2_1sc),
           .msk_a1b0(din_7_msk_ab0), .msk_a1b1(din_7_msk_ab1), .msk_a1b2(din_7_msk_ab2),
           .msk_a1b0_1sc(din_7_msk_ab0_1sc), .msk_a1b1_1sc(din_7_msk_ab1_1sc), .msk_a1b2_1sc(din_7_msk_ab2_1sc),

           .a2b0(din_9_ab0), .a2b1(din_9_ab1),
           .a2b0_1sc(din_9_ab0_1sc), .a2b1_1sc(din_9_ab1_1sc),
           .msk_a2b0(din_9_msk_ab0), .msk_a2b1(din_9_msk_ab1),
           .msk_a2b0_1sc(din_9_msk_ab0_1sc), .msk_a2b1_1sc(din_9_msk_ab1_1sc),
           
           .a3b0(din_11_ab0),
           .a3b0_1sc(din_11_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_6_calc (
           .clk(clk), .sign(din_signs_reg[6]), 
           .p(addr_2_6),
           .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
           .a0b0_1sc(din_6_ab0_1sc), .a0b1_1sc(din_6_ab1_1sc), .a0b2_1sc(din_6_ab2_1sc), .a0b3_1sc(din_6_ab3_1sc),
           .msk_a0b0(din_6_msk_ab0), .msk_a0b1(din_6_msk_ab1), .msk_a0b2(din_6_msk_ab2), .msk_a0b3(din_6_msk_ab3),
           .msk_a0b0_1sc(din_6_msk_ab0_1sc), .msk_a0b1_1sc(din_6_msk_ab1_1sc), .msk_a0b2_1sc(din_6_msk_ab2_1sc), .msk_a0b3_1sc(din_6_msk_ab3_1sc),

           .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2),
           .a1b0_1sc(din_8_ab0_1sc), .a1b1_1sc(din_8_ab1_1sc), .a1b2_1sc(din_8_ab2_1sc),
           .msk_a1b0(din_8_msk_ab0), .msk_a1b1(din_8_msk_ab1), .msk_a1b2(din_8_msk_ab2),
           .msk_a1b0_1sc(din_8_msk_ab0_1sc), .msk_a1b1_1sc(din_8_msk_ab1_1sc), .msk_a1b2_1sc(din_8_msk_ab2_1sc),

           .a2b0(din_10_ab0), .a2b1(din_10_ab1),
           .a2b0_1sc(din_10_ab0_1sc), .a2b1_1sc(din_10_ab1_1sc),
           .msk_a2b0(din_10_msk_ab0), .msk_a2b1(din_10_msk_ab1),
           .msk_a2b0_1sc(din_10_msk_ab0_1sc), .msk_a2b1_1sc(din_10_msk_ab1_1sc),
           
           .a3b0(din_12_ab0),
           .a3b0_1sc(din_12_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_7_calc (
           .clk(clk), .sign(din_signs_reg[7]), 
           .p(addr_2_7),
           .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
           .a0b0_1sc(din_7_ab0_1sc), .a0b1_1sc(din_7_ab1_1sc), .a0b2_1sc(din_7_ab2_1sc), .a0b3_1sc(din_7_ab3_1sc),
           .msk_a0b0(din_7_msk_ab0), .msk_a0b1(din_7_msk_ab1), .msk_a0b2(din_7_msk_ab2), .msk_a0b3(din_7_msk_ab3),
           .msk_a0b0_1sc(din_7_msk_ab0_1sc), .msk_a0b1_1sc(din_7_msk_ab1_1sc), .msk_a0b2_1sc(din_7_msk_ab2_1sc), .msk_a0b3_1sc(din_7_msk_ab3_1sc),

           .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2),
           .a1b0_1sc(din_9_ab0_1sc), .a1b1_1sc(din_9_ab1_1sc), .a1b2_1sc(din_9_ab2_1sc),
           .msk_a1b0(din_9_msk_ab0), .msk_a1b1(din_9_msk_ab1), .msk_a1b2(din_9_msk_ab2),
           .msk_a1b0_1sc(din_9_msk_ab0_1sc), .msk_a1b1_1sc(din_9_msk_ab1_1sc), .msk_a1b2_1sc(din_9_msk_ab2_1sc),

           .a2b0(din_11_ab0), .a2b1(din_11_ab1),
           .a2b0_1sc(din_11_ab0_1sc), .a2b1_1sc(din_11_ab1_1sc),
           .msk_a2b0(din_11_msk_ab0), .msk_a2b1(din_11_msk_ab1),
           .msk_a2b0_1sc(din_11_msk_ab0_1sc), .msk_a2b1_1sc(din_11_msk_ab1_1sc),
           
           .a3b0(din_13_ab0),
           .a3b0_1sc(din_13_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_8_calc (
           .clk(clk), .sign(din_signs_reg[8]), 
           .p(addr_2_8),
           .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
           .a0b0_1sc(din_8_ab0_1sc), .a0b1_1sc(din_8_ab1_1sc), .a0b2_1sc(din_8_ab2_1sc), .a0b3_1sc(din_8_ab3_1sc),
           .msk_a0b0(din_8_msk_ab0), .msk_a0b1(din_8_msk_ab1), .msk_a0b2(din_8_msk_ab2), .msk_a0b3(din_8_msk_ab3),
           .msk_a0b0_1sc(din_8_msk_ab0_1sc), .msk_a0b1_1sc(din_8_msk_ab1_1sc), .msk_a0b2_1sc(din_8_msk_ab2_1sc), .msk_a0b3_1sc(din_8_msk_ab3_1sc),

           .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2),
           .a1b0_1sc(din_10_ab0_1sc), .a1b1_1sc(din_10_ab1_1sc), .a1b2_1sc(din_10_ab2_1sc),
           .msk_a1b0(din_10_msk_ab0), .msk_a1b1(din_10_msk_ab1), .msk_a1b2(din_10_msk_ab2),
           .msk_a1b0_1sc(din_10_msk_ab0_1sc), .msk_a1b1_1sc(din_10_msk_ab1_1sc), .msk_a1b2_1sc(din_10_msk_ab2_1sc),

           .a2b0(din_12_ab0), .a2b1(din_12_ab1),
           .a2b0_1sc(din_12_ab0_1sc), .a2b1_1sc(din_12_ab1_1sc),
           .msk_a2b0(din_12_msk_ab0), .msk_a2b1(din_12_msk_ab1),
           .msk_a2b0_1sc(din_12_msk_ab0_1sc), .msk_a2b1_1sc(din_12_msk_ab1_1sc),
           
           .a3b0(din_14_ab0),
           .a3b0_1sc(din_14_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_9_calc (
           .clk(clk), .sign(din_signs_reg[9]), 
           .p(addr_2_9),
           .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
           .a0b0_1sc(din_9_ab0_1sc), .a0b1_1sc(din_9_ab1_1sc), .a0b2_1sc(din_9_ab2_1sc), .a0b3_1sc(din_9_ab3_1sc),
           .msk_a0b0(din_9_msk_ab0), .msk_a0b1(din_9_msk_ab1), .msk_a0b2(din_9_msk_ab2), .msk_a0b3(din_9_msk_ab3),
           .msk_a0b0_1sc(din_9_msk_ab0_1sc), .msk_a0b1_1sc(din_9_msk_ab1_1sc), .msk_a0b2_1sc(din_9_msk_ab2_1sc), .msk_a0b3_1sc(din_9_msk_ab3_1sc),

           .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2),
           .a1b0_1sc(din_11_ab0_1sc), .a1b1_1sc(din_11_ab1_1sc), .a1b2_1sc(din_11_ab2_1sc),
           .msk_a1b0(din_11_msk_ab0), .msk_a1b1(din_11_msk_ab1), .msk_a1b2(din_11_msk_ab2),
           .msk_a1b0_1sc(din_11_msk_ab0_1sc), .msk_a1b1_1sc(din_11_msk_ab1_1sc), .msk_a1b2_1sc(din_11_msk_ab2_1sc),

           .a2b0(din_13_ab0), .a2b1(din_13_ab1),
           .a2b0_1sc(din_13_ab0_1sc), .a2b1_1sc(din_13_ab1_1sc),
           .msk_a2b0(din_13_msk_ab0), .msk_a2b1(din_13_msk_ab1),
           .msk_a2b0_1sc(din_13_msk_ab0_1sc), .msk_a2b1_1sc(din_13_msk_ab1_1sc),
           
           .a3b0(din_15_ab0),
           .a3b0_1sc(din_15_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_10_calc (
           .clk(clk), .sign(din_signs_reg[10]), 
           .p(addr_2_10),
           .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
           .a0b0_1sc(din_10_ab0_1sc), .a0b1_1sc(din_10_ab1_1sc), .a0b2_1sc(din_10_ab2_1sc), .a0b3_1sc(din_10_ab3_1sc),
           .msk_a0b0(din_10_msk_ab0), .msk_a0b1(din_10_msk_ab1), .msk_a0b2(din_10_msk_ab2), .msk_a0b3(din_10_msk_ab3),
           .msk_a0b0_1sc(din_10_msk_ab0_1sc), .msk_a0b1_1sc(din_10_msk_ab1_1sc), .msk_a0b2_1sc(din_10_msk_ab2_1sc), .msk_a0b3_1sc(din_10_msk_ab3_1sc),

           .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2),
           .a1b0_1sc(din_12_ab0_1sc), .a1b1_1sc(din_12_ab1_1sc), .a1b2_1sc(din_12_ab2_1sc),
           .msk_a1b0(din_12_msk_ab0), .msk_a1b1(din_12_msk_ab1), .msk_a1b2(din_12_msk_ab2),
           .msk_a1b0_1sc(din_12_msk_ab0_1sc), .msk_a1b1_1sc(din_12_msk_ab1_1sc), .msk_a1b2_1sc(din_12_msk_ab2_1sc),

           .a2b0(din_14_ab0), .a2b1(din_14_ab1),
           .a2b0_1sc(din_14_ab0_1sc), .a2b1_1sc(din_14_ab1_1sc),
           .msk_a2b0(din_14_msk_ab0), .msk_a2b1(din_14_msk_ab1),
           .msk_a2b0_1sc(din_14_msk_ab0_1sc), .msk_a2b1_1sc(din_14_msk_ab1_1sc),
           
           .a3b0(din_16_ab0),
           .a3b0_1sc(din_16_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_11_calc (
           .clk(clk), .sign(din_signs_reg[11]), 
           .p(addr_2_11),
           .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
           .a0b0_1sc(din_11_ab0_1sc), .a0b1_1sc(din_11_ab1_1sc), .a0b2_1sc(din_11_ab2_1sc), .a0b3_1sc(din_11_ab3_1sc),
           .msk_a0b0(din_11_msk_ab0), .msk_a0b1(din_11_msk_ab1), .msk_a0b2(din_11_msk_ab2), .msk_a0b3(din_11_msk_ab3),
           .msk_a0b0_1sc(din_11_msk_ab0_1sc), .msk_a0b1_1sc(din_11_msk_ab1_1sc), .msk_a0b2_1sc(din_11_msk_ab2_1sc), .msk_a0b3_1sc(din_11_msk_ab3_1sc),

           .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2),
           .a1b0_1sc(din_13_ab0_1sc), .a1b1_1sc(din_13_ab1_1sc), .a1b2_1sc(din_13_ab2_1sc),
           .msk_a1b0(din_13_msk_ab0), .msk_a1b1(din_13_msk_ab1), .msk_a1b2(din_13_msk_ab2),
           .msk_a1b0_1sc(din_13_msk_ab0_1sc), .msk_a1b1_1sc(din_13_msk_ab1_1sc), .msk_a1b2_1sc(din_13_msk_ab2_1sc),

           .a2b0(din_15_ab0), .a2b1(din_15_ab1),
           .a2b0_1sc(din_15_ab0_1sc), .a2b1_1sc(din_15_ab1_1sc),
           .msk_a2b0(din_15_msk_ab0), .msk_a2b1(din_15_msk_ab1),
           .msk_a2b0_1sc(din_15_msk_ab0_1sc), .msk_a2b1_1sc(din_15_msk_ab1_1sc),
           
           .a3b0(din_17_ab0),
           .a3b0_1sc(din_17_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_12_calc (
           .clk(clk), .sign(din_signs_reg[12]), 
           .p(addr_2_12),
           .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
           .a0b0_1sc(din_12_ab0_1sc), .a0b1_1sc(din_12_ab1_1sc), .a0b2_1sc(din_12_ab2_1sc), .a0b3_1sc(din_12_ab3_1sc),
           .msk_a0b0(din_12_msk_ab0), .msk_a0b1(din_12_msk_ab1), .msk_a0b2(din_12_msk_ab2), .msk_a0b3(din_12_msk_ab3),
           .msk_a0b0_1sc(din_12_msk_ab0_1sc), .msk_a0b1_1sc(din_12_msk_ab1_1sc), .msk_a0b2_1sc(din_12_msk_ab2_1sc), .msk_a0b3_1sc(din_12_msk_ab3_1sc),

           .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2),
           .a1b0_1sc(din_14_ab0_1sc), .a1b1_1sc(din_14_ab1_1sc), .a1b2_1sc(din_14_ab2_1sc),
           .msk_a1b0(din_14_msk_ab0), .msk_a1b1(din_14_msk_ab1), .msk_a1b2(din_14_msk_ab2),
           .msk_a1b0_1sc(din_14_msk_ab0_1sc), .msk_a1b1_1sc(din_14_msk_ab1_1sc), .msk_a1b2_1sc(din_14_msk_ab2_1sc),

           .a2b0(din_16_ab0), .a2b1(din_16_ab1),
           .a2b0_1sc(din_16_ab0_1sc), .a2b1_1sc(din_16_ab1_1sc),
           .msk_a2b0(din_16_msk_ab0), .msk_a2b1(din_16_msk_ab1),
           .msk_a2b0_1sc(din_16_msk_ab0_1sc), .msk_a2b1_1sc(din_16_msk_ab1_1sc),
           
           .a3b0(din_18_ab0),
           .a3b0_1sc(din_18_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_13_calc (
           .clk(clk), .sign(din_signs_reg[13]), 
           .p(addr_2_13),
           .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
           .a0b0_1sc(din_13_ab0_1sc), .a0b1_1sc(din_13_ab1_1sc), .a0b2_1sc(din_13_ab2_1sc), .a0b3_1sc(din_13_ab3_1sc),
           .msk_a0b0(din_13_msk_ab0), .msk_a0b1(din_13_msk_ab1), .msk_a0b2(din_13_msk_ab2), .msk_a0b3(din_13_msk_ab3),
           .msk_a0b0_1sc(din_13_msk_ab0_1sc), .msk_a0b1_1sc(din_13_msk_ab1_1sc), .msk_a0b2_1sc(din_13_msk_ab2_1sc), .msk_a0b3_1sc(din_13_msk_ab3_1sc),

           .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2),
           .a1b0_1sc(din_15_ab0_1sc), .a1b1_1sc(din_15_ab1_1sc), .a1b2_1sc(din_15_ab2_1sc),
           .msk_a1b0(din_15_msk_ab0), .msk_a1b1(din_15_msk_ab1), .msk_a1b2(din_15_msk_ab2),
           .msk_a1b0_1sc(din_15_msk_ab0_1sc), .msk_a1b1_1sc(din_15_msk_ab1_1sc), .msk_a1b2_1sc(din_15_msk_ab2_1sc),

           .a2b0(din_17_ab0), .a2b1(din_17_ab1),
           .a2b0_1sc(din_17_ab0_1sc), .a2b1_1sc(din_17_ab1_1sc),
           .msk_a2b0(din_17_msk_ab0), .msk_a2b1(din_17_msk_ab1),
           .msk_a2b0_1sc(din_17_msk_ab0_1sc), .msk_a2b1_1sc(din_17_msk_ab1_1sc),
           
           .a3b0(din_19_ab0),
           .a3b0_1sc(din_19_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_14_calc (
           .clk(clk), .sign(din_signs_reg[14]), 
           .p(addr_2_14),
           .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
           .a0b0_1sc(din_14_ab0_1sc), .a0b1_1sc(din_14_ab1_1sc), .a0b2_1sc(din_14_ab2_1sc), .a0b3_1sc(din_14_ab3_1sc),
           .msk_a0b0(din_14_msk_ab0), .msk_a0b1(din_14_msk_ab1), .msk_a0b2(din_14_msk_ab2), .msk_a0b3(din_14_msk_ab3),
           .msk_a0b0_1sc(din_14_msk_ab0_1sc), .msk_a0b1_1sc(din_14_msk_ab1_1sc), .msk_a0b2_1sc(din_14_msk_ab2_1sc), .msk_a0b3_1sc(din_14_msk_ab3_1sc),

           .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2),
           .a1b0_1sc(din_16_ab0_1sc), .a1b1_1sc(din_16_ab1_1sc), .a1b2_1sc(din_16_ab2_1sc),
           .msk_a1b0(din_16_msk_ab0), .msk_a1b1(din_16_msk_ab1), .msk_a1b2(din_16_msk_ab2),
           .msk_a1b0_1sc(din_16_msk_ab0_1sc), .msk_a1b1_1sc(din_16_msk_ab1_1sc), .msk_a1b2_1sc(din_16_msk_ab2_1sc),

           .a2b0(din_18_ab0), .a2b1(din_18_ab1),
           .a2b0_1sc(din_18_ab0_1sc), .a2b1_1sc(din_18_ab1_1sc),
           .msk_a2b0(din_18_msk_ab0), .msk_a2b1(din_18_msk_ab1),
           .msk_a2b0_1sc(din_18_msk_ab0_1sc), .msk_a2b1_1sc(din_18_msk_ab1_1sc),
           
           .a3b0(din_20_ab0),
           .a3b0_1sc(din_20_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_15_calc (
           .clk(clk), .sign(din_signs_reg[15]), 
           .p(addr_2_15),
           .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
           .a0b0_1sc(din_15_ab0_1sc), .a0b1_1sc(din_15_ab1_1sc), .a0b2_1sc(din_15_ab2_1sc), .a0b3_1sc(din_15_ab3_1sc),
           .msk_a0b0(din_15_msk_ab0), .msk_a0b1(din_15_msk_ab1), .msk_a0b2(din_15_msk_ab2), .msk_a0b3(din_15_msk_ab3),
           .msk_a0b0_1sc(din_15_msk_ab0_1sc), .msk_a0b1_1sc(din_15_msk_ab1_1sc), .msk_a0b2_1sc(din_15_msk_ab2_1sc), .msk_a0b3_1sc(din_15_msk_ab3_1sc),

           .a1b0(din_17_ab0), .a1b1(din_17_ab1), .a1b2(din_17_ab2),
           .a1b0_1sc(din_17_ab0_1sc), .a1b1_1sc(din_17_ab1_1sc), .a1b2_1sc(din_17_ab2_1sc),
           .msk_a1b0(din_17_msk_ab0), .msk_a1b1(din_17_msk_ab1), .msk_a1b2(din_17_msk_ab2),
           .msk_a1b0_1sc(din_17_msk_ab0_1sc), .msk_a1b1_1sc(din_17_msk_ab1_1sc), .msk_a1b2_1sc(din_17_msk_ab2_1sc),

           .a2b0(din_19_ab0), .a2b1(din_19_ab1),
           .a2b0_1sc(din_19_ab0_1sc), .a2b1_1sc(din_19_ab1_1sc),
           .msk_a2b0(din_19_msk_ab0), .msk_a2b1(din_19_msk_ab1),
           .msk_a2b0_1sc(din_19_msk_ab0_1sc), .msk_a2b1_1sc(din_19_msk_ab1_1sc),
           
           .a3b0(din_21_ab0),
           .a3b0_1sc(din_21_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_16_calc (
           .clk(clk), .sign(din_signs_reg[16]), 
           .p(addr_2_16),
           .a0b0(din_16_ab0), .a0b1(din_16_ab1), .a0b2(din_16_ab2), .a0b3(din_16_ab3),
           .a0b0_1sc(din_16_ab0_1sc), .a0b1_1sc(din_16_ab1_1sc), .a0b2_1sc(din_16_ab2_1sc), .a0b3_1sc(din_16_ab3_1sc),
           .msk_a0b0(din_16_msk_ab0), .msk_a0b1(din_16_msk_ab1), .msk_a0b2(din_16_msk_ab2), .msk_a0b3(din_16_msk_ab3),
           .msk_a0b0_1sc(din_16_msk_ab0_1sc), .msk_a0b1_1sc(din_16_msk_ab1_1sc), .msk_a0b2_1sc(din_16_msk_ab2_1sc), .msk_a0b3_1sc(din_16_msk_ab3_1sc),

           .a1b0(din_18_ab0), .a1b1(din_18_ab1), .a1b2(din_18_ab2),
           .a1b0_1sc(din_18_ab0_1sc), .a1b1_1sc(din_18_ab1_1sc), .a1b2_1sc(din_18_ab2_1sc),
           .msk_a1b0(din_18_msk_ab0), .msk_a1b1(din_18_msk_ab1), .msk_a1b2(din_18_msk_ab2),
           .msk_a1b0_1sc(din_18_msk_ab0_1sc), .msk_a1b1_1sc(din_18_msk_ab1_1sc), .msk_a1b2_1sc(din_18_msk_ab2_1sc),

           .a2b0(din_20_ab0), .a2b1(din_20_ab1),
           .a2b0_1sc(din_20_ab0_1sc), .a2b1_1sc(din_20_ab1_1sc),
           .msk_a2b0(din_20_msk_ab0), .msk_a2b1(din_20_msk_ab1),
           .msk_a2b0_1sc(din_20_msk_ab0_1sc), .msk_a2b1_1sc(din_20_msk_ab1_1sc),
           
           .a3b0(din_22_ab0),
           .a3b0_1sc(din_22_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_17_calc (
           .clk(clk), .sign(din_signs_reg[17]), 
           .p(addr_2_17),
           .a0b0(din_17_ab0), .a0b1(din_17_ab1), .a0b2(din_17_ab2), .a0b3(din_17_ab3),
           .a0b0_1sc(din_17_ab0_1sc), .a0b1_1sc(din_17_ab1_1sc), .a0b2_1sc(din_17_ab2_1sc), .a0b3_1sc(din_17_ab3_1sc),
           .msk_a0b0(din_17_msk_ab0), .msk_a0b1(din_17_msk_ab1), .msk_a0b2(din_17_msk_ab2), .msk_a0b3(din_17_msk_ab3),
           .msk_a0b0_1sc(din_17_msk_ab0_1sc), .msk_a0b1_1sc(din_17_msk_ab1_1sc), .msk_a0b2_1sc(din_17_msk_ab2_1sc), .msk_a0b3_1sc(din_17_msk_ab3_1sc),

           .a1b0(din_19_ab0), .a1b1(din_19_ab1), .a1b2(din_19_ab2),
           .a1b0_1sc(din_19_ab0_1sc), .a1b1_1sc(din_19_ab1_1sc), .a1b2_1sc(din_19_ab2_1sc),
           .msk_a1b0(din_19_msk_ab0), .msk_a1b1(din_19_msk_ab1), .msk_a1b2(din_19_msk_ab2),
           .msk_a1b0_1sc(din_19_msk_ab0_1sc), .msk_a1b1_1sc(din_19_msk_ab1_1sc), .msk_a1b2_1sc(din_19_msk_ab2_1sc),

           .a2b0(din_21_ab0), .a2b1(din_21_ab1),
           .a2b0_1sc(din_21_ab0_1sc), .a2b1_1sc(din_21_ab1_1sc),
           .msk_a2b0(din_21_msk_ab0), .msk_a2b1(din_21_msk_ab1),
           .msk_a2b0_1sc(din_21_msk_ab0_1sc), .msk_a2b1_1sc(din_21_msk_ab1_1sc),
           
           .a3b0(din_23_ab0),
           .a3b0_1sc(din_23_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_18_calc (
           .clk(clk), .sign(din_signs_reg[18]), 
           .p(addr_2_18),
           .a0b0(din_18_ab0), .a0b1(din_18_ab1), .a0b2(din_18_ab2), .a0b3(din_18_ab3),
           .a0b0_1sc(din_18_ab0_1sc), .a0b1_1sc(din_18_ab1_1sc), .a0b2_1sc(din_18_ab2_1sc), .a0b3_1sc(din_18_ab3_1sc),
           .msk_a0b0(din_18_msk_ab0), .msk_a0b1(din_18_msk_ab1), .msk_a0b2(din_18_msk_ab2), .msk_a0b3(din_18_msk_ab3),
           .msk_a0b0_1sc(din_18_msk_ab0_1sc), .msk_a0b1_1sc(din_18_msk_ab1_1sc), .msk_a0b2_1sc(din_18_msk_ab2_1sc), .msk_a0b3_1sc(din_18_msk_ab3_1sc),

           .a1b0(din_20_ab0), .a1b1(din_20_ab1), .a1b2(din_20_ab2),
           .a1b0_1sc(din_20_ab0_1sc), .a1b1_1sc(din_20_ab1_1sc), .a1b2_1sc(din_20_ab2_1sc),
           .msk_a1b0(din_20_msk_ab0), .msk_a1b1(din_20_msk_ab1), .msk_a1b2(din_20_msk_ab2),
           .msk_a1b0_1sc(din_20_msk_ab0_1sc), .msk_a1b1_1sc(din_20_msk_ab1_1sc), .msk_a1b2_1sc(din_20_msk_ab2_1sc),

           .a2b0(din_22_ab0), .a2b1(din_22_ab1),
           .a2b0_1sc(din_22_ab0_1sc), .a2b1_1sc(din_22_ab1_1sc),
           .msk_a2b0(din_22_msk_ab0), .msk_a2b1(din_22_msk_ab1),
           .msk_a2b0_1sc(din_22_msk_ab0_1sc), .msk_a2b1_1sc(din_22_msk_ab1_1sc),
           
           .a3b0(din_24_ab0),
           .a3b0_1sc(din_24_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_19_calc (
           .clk(clk), .sign(din_signs_reg[19]), 
           .p(addr_2_19),
           .a0b0(din_19_ab0), .a0b1(din_19_ab1), .a0b2(din_19_ab2), .a0b3(din_19_ab3),
           .a0b0_1sc(din_19_ab0_1sc), .a0b1_1sc(din_19_ab1_1sc), .a0b2_1sc(din_19_ab2_1sc), .a0b3_1sc(din_19_ab3_1sc),
           .msk_a0b0(din_19_msk_ab0), .msk_a0b1(din_19_msk_ab1), .msk_a0b2(din_19_msk_ab2), .msk_a0b3(din_19_msk_ab3),
           .msk_a0b0_1sc(din_19_msk_ab0_1sc), .msk_a0b1_1sc(din_19_msk_ab1_1sc), .msk_a0b2_1sc(din_19_msk_ab2_1sc), .msk_a0b3_1sc(din_19_msk_ab3_1sc),

           .a1b0(din_21_ab0), .a1b1(din_21_ab1), .a1b2(din_21_ab2),
           .a1b0_1sc(din_21_ab0_1sc), .a1b1_1sc(din_21_ab1_1sc), .a1b2_1sc(din_21_ab2_1sc),
           .msk_a1b0(din_21_msk_ab0), .msk_a1b1(din_21_msk_ab1), .msk_a1b2(din_21_msk_ab2),
           .msk_a1b0_1sc(din_21_msk_ab0_1sc), .msk_a1b1_1sc(din_21_msk_ab1_1sc), .msk_a1b2_1sc(din_21_msk_ab2_1sc),

           .a2b0(din_23_ab0), .a2b1(din_23_ab1),
           .a2b0_1sc(din_23_ab0_1sc), .a2b1_1sc(din_23_ab1_1sc),
           .msk_a2b0(din_23_msk_ab0), .msk_a2b1(din_23_msk_ab1),
           .msk_a2b0_1sc(din_23_msk_ab0_1sc), .msk_a2b1_1sc(din_23_msk_ab1_1sc),
           
           .a3b0(din_25_ab0),
           .a3b0_1sc(din_25_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_20_calc (
           .clk(clk), .sign(din_signs_reg[20]), 
           .p(addr_2_20),
           .a0b0(din_20_ab0), .a0b1(din_20_ab1), .a0b2(din_20_ab2), .a0b3(din_20_ab3),
           .a0b0_1sc(din_20_ab0_1sc), .a0b1_1sc(din_20_ab1_1sc), .a0b2_1sc(din_20_ab2_1sc), .a0b3_1sc(din_20_ab3_1sc),
           .msk_a0b0(din_20_msk_ab0), .msk_a0b1(din_20_msk_ab1), .msk_a0b2(din_20_msk_ab2), .msk_a0b3(din_20_msk_ab3),
           .msk_a0b0_1sc(din_20_msk_ab0_1sc), .msk_a0b1_1sc(din_20_msk_ab1_1sc), .msk_a0b2_1sc(din_20_msk_ab2_1sc), .msk_a0b3_1sc(din_20_msk_ab3_1sc),

           .a1b0(din_22_ab0), .a1b1(din_22_ab1), .a1b2(din_22_ab2),
           .a1b0_1sc(din_22_ab0_1sc), .a1b1_1sc(din_22_ab1_1sc), .a1b2_1sc(din_22_ab2_1sc),
           .msk_a1b0(din_22_msk_ab0), .msk_a1b1(din_22_msk_ab1), .msk_a1b2(din_22_msk_ab2),
           .msk_a1b0_1sc(din_22_msk_ab0_1sc), .msk_a1b1_1sc(din_22_msk_ab1_1sc), .msk_a1b2_1sc(din_22_msk_ab2_1sc),

           .a2b0(din_24_ab0), .a2b1(din_24_ab1),
           .a2b0_1sc(din_24_ab0_1sc), .a2b1_1sc(din_24_ab1_1sc),
           .msk_a2b0(din_24_msk_ab0), .msk_a2b1(din_24_msk_ab1),
           .msk_a2b0_1sc(din_24_msk_ab0_1sc), .msk_a2b1_1sc(din_24_msk_ab1_1sc),
           
           .a3b0(din_26_ab0),
           .a3b0_1sc(din_26_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_21_calc (
           .clk(clk), .sign(din_signs_reg[21]), 
           .p(addr_2_21),
           .a0b0(din_21_ab0), .a0b1(din_21_ab1), .a0b2(din_21_ab2), .a0b3(din_21_ab3),
           .a0b0_1sc(din_21_ab0_1sc), .a0b1_1sc(din_21_ab1_1sc), .a0b2_1sc(din_21_ab2_1sc), .a0b3_1sc(din_21_ab3_1sc),
           .msk_a0b0(din_21_msk_ab0), .msk_a0b1(din_21_msk_ab1), .msk_a0b2(din_21_msk_ab2), .msk_a0b3(din_21_msk_ab3),
           .msk_a0b0_1sc(din_21_msk_ab0_1sc), .msk_a0b1_1sc(din_21_msk_ab1_1sc), .msk_a0b2_1sc(din_21_msk_ab2_1sc), .msk_a0b3_1sc(din_21_msk_ab3_1sc),

           .a1b0(din_23_ab0), .a1b1(din_23_ab1), .a1b2(din_23_ab2),
           .a1b0_1sc(din_23_ab0_1sc), .a1b1_1sc(din_23_ab1_1sc), .a1b2_1sc(din_23_ab2_1sc),
           .msk_a1b0(din_23_msk_ab0), .msk_a1b1(din_23_msk_ab1), .msk_a1b2(din_23_msk_ab2),
           .msk_a1b0_1sc(din_23_msk_ab0_1sc), .msk_a1b1_1sc(din_23_msk_ab1_1sc), .msk_a1b2_1sc(din_23_msk_ab2_1sc),

           .a2b0(din_25_ab0), .a2b1(din_25_ab1),
           .a2b0_1sc(din_25_ab0_1sc), .a2b1_1sc(din_25_ab1_1sc),
           .msk_a2b0(din_25_msk_ab0), .msk_a2b1(din_25_msk_ab1),
           .msk_a2b0_1sc(din_25_msk_ab0_1sc), .msk_a2b1_1sc(din_25_msk_ab1_1sc),
           
           .a3b0(din_27_ab0),
           .a3b0_1sc(din_27_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_22_calc (
           .clk(clk), .sign(din_signs_reg[22]), 
           .p(addr_2_22),
           .a0b0(din_22_ab0), .a0b1(din_22_ab1), .a0b2(din_22_ab2), .a0b3(din_22_ab3),
           .a0b0_1sc(din_22_ab0_1sc), .a0b1_1sc(din_22_ab1_1sc), .a0b2_1sc(din_22_ab2_1sc), .a0b3_1sc(din_22_ab3_1sc),
           .msk_a0b0(din_22_msk_ab0), .msk_a0b1(din_22_msk_ab1), .msk_a0b2(din_22_msk_ab2), .msk_a0b3(din_22_msk_ab3),
           .msk_a0b0_1sc(din_22_msk_ab0_1sc), .msk_a0b1_1sc(din_22_msk_ab1_1sc), .msk_a0b2_1sc(din_22_msk_ab2_1sc), .msk_a0b3_1sc(din_22_msk_ab3_1sc),

           .a1b0(din_24_ab0), .a1b1(din_24_ab1), .a1b2(din_24_ab2),
           .a1b0_1sc(din_24_ab0_1sc), .a1b1_1sc(din_24_ab1_1sc), .a1b2_1sc(din_24_ab2_1sc),
           .msk_a1b0(din_24_msk_ab0), .msk_a1b1(din_24_msk_ab1), .msk_a1b2(din_24_msk_ab2),
           .msk_a1b0_1sc(din_24_msk_ab0_1sc), .msk_a1b1_1sc(din_24_msk_ab1_1sc), .msk_a1b2_1sc(din_24_msk_ab2_1sc),

           .a2b0(din_26_ab0), .a2b1(din_26_ab1),
           .a2b0_1sc(din_26_ab0_1sc), .a2b1_1sc(din_26_ab1_1sc),
           .msk_a2b0(din_26_msk_ab0), .msk_a2b1(din_26_msk_ab1),
           .msk_a2b0_1sc(din_26_msk_ab0_1sc), .msk_a2b1_1sc(din_26_msk_ab1_1sc),
           
           .a3b0(din_28_ab0),
           .a3b0_1sc(din_28_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_23_calc (
           .clk(clk), .sign(din_signs_reg[23]), 
           .p(addr_2_23),
           .a0b0(din_23_ab0), .a0b1(din_23_ab1), .a0b2(din_23_ab2), .a0b3(din_23_ab3),
           .a0b0_1sc(din_23_ab0_1sc), .a0b1_1sc(din_23_ab1_1sc), .a0b2_1sc(din_23_ab2_1sc), .a0b3_1sc(din_23_ab3_1sc),
           .msk_a0b0(din_23_msk_ab0), .msk_a0b1(din_23_msk_ab1), .msk_a0b2(din_23_msk_ab2), .msk_a0b3(din_23_msk_ab3),
           .msk_a0b0_1sc(din_23_msk_ab0_1sc), .msk_a0b1_1sc(din_23_msk_ab1_1sc), .msk_a0b2_1sc(din_23_msk_ab2_1sc), .msk_a0b3_1sc(din_23_msk_ab3_1sc),

           .a1b0(din_25_ab0), .a1b1(din_25_ab1), .a1b2(din_25_ab2),
           .a1b0_1sc(din_25_ab0_1sc), .a1b1_1sc(din_25_ab1_1sc), .a1b2_1sc(din_25_ab2_1sc),
           .msk_a1b0(din_25_msk_ab0), .msk_a1b1(din_25_msk_ab1), .msk_a1b2(din_25_msk_ab2),
           .msk_a1b0_1sc(din_25_msk_ab0_1sc), .msk_a1b1_1sc(din_25_msk_ab1_1sc), .msk_a1b2_1sc(din_25_msk_ab2_1sc),

           .a2b0(din_27_ab0), .a2b1(din_27_ab1),
           .a2b0_1sc(din_27_ab0_1sc), .a2b1_1sc(din_27_ab1_1sc),
           .msk_a2b0(din_27_msk_ab0), .msk_a2b1(din_27_msk_ab1),
           .msk_a2b0_1sc(din_27_msk_ab0_1sc), .msk_a2b1_1sc(din_27_msk_ab1_1sc),
           
           .a3b0(din_29_ab0),
           .a3b0_1sc(din_29_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_24_calc (
           .clk(clk), .sign(din_signs_reg[24]), 
           .p(addr_2_24),
           .a0b0(din_24_ab0), .a0b1(din_24_ab1), .a0b2(din_24_ab2), .a0b3(din_24_ab3),
           .a0b0_1sc(din_24_ab0_1sc), .a0b1_1sc(din_24_ab1_1sc), .a0b2_1sc(din_24_ab2_1sc), .a0b3_1sc(din_24_ab3_1sc),
           .msk_a0b0(din_24_msk_ab0), .msk_a0b1(din_24_msk_ab1), .msk_a0b2(din_24_msk_ab2), .msk_a0b3(din_24_msk_ab3),
           .msk_a0b0_1sc(din_24_msk_ab0_1sc), .msk_a0b1_1sc(din_24_msk_ab1_1sc), .msk_a0b2_1sc(din_24_msk_ab2_1sc), .msk_a0b3_1sc(din_24_msk_ab3_1sc),

           .a1b0(din_26_ab0), .a1b1(din_26_ab1), .a1b2(din_26_ab2),
           .a1b0_1sc(din_26_ab0_1sc), .a1b1_1sc(din_26_ab1_1sc), .a1b2_1sc(din_26_ab2_1sc),
           .msk_a1b0(din_26_msk_ab0), .msk_a1b1(din_26_msk_ab1), .msk_a1b2(din_26_msk_ab2),
           .msk_a1b0_1sc(din_26_msk_ab0_1sc), .msk_a1b1_1sc(din_26_msk_ab1_1sc), .msk_a1b2_1sc(din_26_msk_ab2_1sc),

           .a2b0(din_28_ab0), .a2b1(din_28_ab1),
           .a2b0_1sc(din_28_ab0_1sc), .a2b1_1sc(din_28_ab1_1sc),
           .msk_a2b0(din_28_msk_ab0), .msk_a2b1(din_28_msk_ab1),
           .msk_a2b0_1sc(din_28_msk_ab0_1sc), .msk_a2b1_1sc(din_28_msk_ab1_1sc),
           
           .a3b0(din_30_ab0),
           .a3b0_1sc(din_30_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_25_calc (
           .clk(clk), .sign(din_signs_reg[25]), 
           .p(addr_2_25),
           .a0b0(din_25_ab0), .a0b1(din_25_ab1), .a0b2(din_25_ab2), .a0b3(din_25_ab3),
           .a0b0_1sc(din_25_ab0_1sc), .a0b1_1sc(din_25_ab1_1sc), .a0b2_1sc(din_25_ab2_1sc), .a0b3_1sc(din_25_ab3_1sc),
           .msk_a0b0(din_25_msk_ab0), .msk_a0b1(din_25_msk_ab1), .msk_a0b2(din_25_msk_ab2), .msk_a0b3(din_25_msk_ab3),
           .msk_a0b0_1sc(din_25_msk_ab0_1sc), .msk_a0b1_1sc(din_25_msk_ab1_1sc), .msk_a0b2_1sc(din_25_msk_ab2_1sc), .msk_a0b3_1sc(din_25_msk_ab3_1sc),

           .a1b0(din_27_ab0), .a1b1(din_27_ab1), .a1b2(din_27_ab2),
           .a1b0_1sc(din_27_ab0_1sc), .a1b1_1sc(din_27_ab1_1sc), .a1b2_1sc(din_27_ab2_1sc),
           .msk_a1b0(din_27_msk_ab0), .msk_a1b1(din_27_msk_ab1), .msk_a1b2(din_27_msk_ab2),
           .msk_a1b0_1sc(din_27_msk_ab0_1sc), .msk_a1b1_1sc(din_27_msk_ab1_1sc), .msk_a1b2_1sc(din_27_msk_ab2_1sc),

           .a2b0(din_29_ab0), .a2b1(din_29_ab1),
           .a2b0_1sc(din_29_ab0_1sc), .a2b1_1sc(din_29_ab1_1sc),
           .msk_a2b0(din_29_msk_ab0), .msk_a2b1(din_29_msk_ab1),
           .msk_a2b0_1sc(din_29_msk_ab0_1sc), .msk_a2b1_1sc(din_29_msk_ab1_1sc),
           
           .a3b0(din_31_ab0),
           .a3b0_1sc(din_31_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_26_calc (
           .clk(clk), .sign(din_signs_reg[26]), 
           .p(addr_2_26),
           .a0b0(din_26_ab0), .a0b1(din_26_ab1), .a0b2(din_26_ab2), .a0b3(din_26_ab3),
           .a0b0_1sc(din_26_ab0_1sc), .a0b1_1sc(din_26_ab1_1sc), .a0b2_1sc(din_26_ab2_1sc), .a0b3_1sc(din_26_ab3_1sc),
           .msk_a0b0(din_26_msk_ab0), .msk_a0b1(din_26_msk_ab1), .msk_a0b2(din_26_msk_ab2), .msk_a0b3(din_26_msk_ab3),
           .msk_a0b0_1sc(din_26_msk_ab0_1sc), .msk_a0b1_1sc(din_26_msk_ab1_1sc), .msk_a0b2_1sc(din_26_msk_ab2_1sc), .msk_a0b3_1sc(din_26_msk_ab3_1sc),

           .a1b0(din_28_ab0), .a1b1(din_28_ab1), .a1b2(din_28_ab2),
           .a1b0_1sc(din_28_ab0_1sc), .a1b1_1sc(din_28_ab1_1sc), .a1b2_1sc(din_28_ab2_1sc),
           .msk_a1b0(din_28_msk_ab0), .msk_a1b1(din_28_msk_ab1), .msk_a1b2(din_28_msk_ab2),
           .msk_a1b0_1sc(din_28_msk_ab0_1sc), .msk_a1b1_1sc(din_28_msk_ab1_1sc), .msk_a1b2_1sc(din_28_msk_ab2_1sc),

           .a2b0(din_30_ab0), .a2b1(din_30_ab1),
           .a2b0_1sc(din_30_ab0_1sc), .a2b1_1sc(din_30_ab1_1sc),
           .msk_a2b0(din_30_msk_ab0), .msk_a2b1(din_30_msk_ab1),
           .msk_a2b0_1sc(din_30_msk_ab0_1sc), .msk_a2b1_1sc(din_30_msk_ab1_1sc),
           
           .a3b0(din_32_ab0),
           .a3b0_1sc(din_32_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_27_calc (
           .clk(clk), .sign(din_signs_reg[27]), 
           .p(addr_2_27),
           .a0b0(din_27_ab0), .a0b1(din_27_ab1), .a0b2(din_27_ab2), .a0b3(din_27_ab3),
           .a0b0_1sc(din_27_ab0_1sc), .a0b1_1sc(din_27_ab1_1sc), .a0b2_1sc(din_27_ab2_1sc), .a0b3_1sc(din_27_ab3_1sc),
           .msk_a0b0(din_27_msk_ab0), .msk_a0b1(din_27_msk_ab1), .msk_a0b2(din_27_msk_ab2), .msk_a0b3(din_27_msk_ab3),
           .msk_a0b0_1sc(din_27_msk_ab0_1sc), .msk_a0b1_1sc(din_27_msk_ab1_1sc), .msk_a0b2_1sc(din_27_msk_ab2_1sc), .msk_a0b3_1sc(din_27_msk_ab3_1sc),

           .a1b0(din_29_ab0), .a1b1(din_29_ab1), .a1b2(din_29_ab2),
           .a1b0_1sc(din_29_ab0_1sc), .a1b1_1sc(din_29_ab1_1sc), .a1b2_1sc(din_29_ab2_1sc),
           .msk_a1b0(din_29_msk_ab0), .msk_a1b1(din_29_msk_ab1), .msk_a1b2(din_29_msk_ab2),
           .msk_a1b0_1sc(din_29_msk_ab0_1sc), .msk_a1b1_1sc(din_29_msk_ab1_1sc), .msk_a1b2_1sc(din_29_msk_ab2_1sc),

           .a2b0(din_31_ab0), .a2b1(din_31_ab1),
           .a2b0_1sc(din_31_ab0_1sc), .a2b1_1sc(din_31_ab1_1sc),
           .msk_a2b0(din_31_msk_ab0), .msk_a2b1(din_31_msk_ab1),
           .msk_a2b0_1sc(din_31_msk_ab0_1sc), .msk_a2b1_1sc(din_31_msk_ab1_1sc),
           
           .a3b0(din_33_ab0),
           .a3b0_1sc(din_33_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_28_calc (
           .clk(clk), .sign(din_signs_reg[28]), 
           .p(addr_2_28),
           .a0b0(din_28_ab0), .a0b1(din_28_ab1), .a0b2(din_28_ab2), .a0b3(din_28_ab3),
           .a0b0_1sc(din_28_ab0_1sc), .a0b1_1sc(din_28_ab1_1sc), .a0b2_1sc(din_28_ab2_1sc), .a0b3_1sc(din_28_ab3_1sc),
           .msk_a0b0(din_28_msk_ab0), .msk_a0b1(din_28_msk_ab1), .msk_a0b2(din_28_msk_ab2), .msk_a0b3(din_28_msk_ab3),
           .msk_a0b0_1sc(din_28_msk_ab0_1sc), .msk_a0b1_1sc(din_28_msk_ab1_1sc), .msk_a0b2_1sc(din_28_msk_ab2_1sc), .msk_a0b3_1sc(din_28_msk_ab3_1sc),

           .a1b0(din_30_ab0), .a1b1(din_30_ab1), .a1b2(din_30_ab2),
           .a1b0_1sc(din_30_ab0_1sc), .a1b1_1sc(din_30_ab1_1sc), .a1b2_1sc(din_30_ab2_1sc),
           .msk_a1b0(din_30_msk_ab0), .msk_a1b1(din_30_msk_ab1), .msk_a1b2(din_30_msk_ab2),
           .msk_a1b0_1sc(din_30_msk_ab0_1sc), .msk_a1b1_1sc(din_30_msk_ab1_1sc), .msk_a1b2_1sc(din_30_msk_ab2_1sc),

           .a2b0(din_32_ab0), .a2b1(din_32_ab1),
           .a2b0_1sc(din_32_ab0_1sc), .a2b1_1sc(din_32_ab1_1sc),
           .msk_a2b0(din_32_msk_ab0), .msk_a2b1(din_32_msk_ab1),
           .msk_a2b0_1sc(din_32_msk_ab0_1sc), .msk_a2b1_1sc(din_32_msk_ab1_1sc),
           
           .a3b0(din_34_ab0),
           .a3b0_1sc(din_34_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_29_calc (
           .clk(clk), .sign(din_signs_reg[29]), 
           .p(addr_2_29),
           .a0b0(din_29_ab0), .a0b1(din_29_ab1), .a0b2(din_29_ab2), .a0b3(din_29_ab3),
           .a0b0_1sc(din_29_ab0_1sc), .a0b1_1sc(din_29_ab1_1sc), .a0b2_1sc(din_29_ab2_1sc), .a0b3_1sc(din_29_ab3_1sc),
           .msk_a0b0(din_29_msk_ab0), .msk_a0b1(din_29_msk_ab1), .msk_a0b2(din_29_msk_ab2), .msk_a0b3(din_29_msk_ab3),
           .msk_a0b0_1sc(din_29_msk_ab0_1sc), .msk_a0b1_1sc(din_29_msk_ab1_1sc), .msk_a0b2_1sc(din_29_msk_ab2_1sc), .msk_a0b3_1sc(din_29_msk_ab3_1sc),

           .a1b0(din_31_ab0), .a1b1(din_31_ab1), .a1b2(din_31_ab2),
           .a1b0_1sc(din_31_ab0_1sc), .a1b1_1sc(din_31_ab1_1sc), .a1b2_1sc(din_31_ab2_1sc),
           .msk_a1b0(din_31_msk_ab0), .msk_a1b1(din_31_msk_ab1), .msk_a1b2(din_31_msk_ab2),
           .msk_a1b0_1sc(din_31_msk_ab0_1sc), .msk_a1b1_1sc(din_31_msk_ab1_1sc), .msk_a1b2_1sc(din_31_msk_ab2_1sc),

           .a2b0(din_33_ab0), .a2b1(din_33_ab1),
           .a2b0_1sc(din_33_ab0_1sc), .a2b1_1sc(din_33_ab1_1sc),
           .msk_a2b0(din_33_msk_ab0), .msk_a2b1(din_33_msk_ab1),
           .msk_a2b0_1sc(din_33_msk_ab0_1sc), .msk_a2b1_1sc(din_33_msk_ab1_1sc),
           
           .a3b0(din_35_ab0),
           .a3b0_1sc(din_35_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_30_calc (
           .clk(clk), .sign(din_signs_reg[30]), 
           .p(addr_2_30),
           .a0b0(din_30_ab0), .a0b1(din_30_ab1), .a0b2(din_30_ab2), .a0b3(din_30_ab3),
           .a0b0_1sc(din_30_ab0_1sc), .a0b1_1sc(din_30_ab1_1sc), .a0b2_1sc(din_30_ab2_1sc), .a0b3_1sc(din_30_ab3_1sc),
           .msk_a0b0(din_30_msk_ab0), .msk_a0b1(din_30_msk_ab1), .msk_a0b2(din_30_msk_ab2), .msk_a0b3(din_30_msk_ab3),
           .msk_a0b0_1sc(din_30_msk_ab0_1sc), .msk_a0b1_1sc(din_30_msk_ab1_1sc), .msk_a0b2_1sc(din_30_msk_ab2_1sc), .msk_a0b3_1sc(din_30_msk_ab3_1sc),

           .a1b0(din_32_ab0), .a1b1(din_32_ab1), .a1b2(din_32_ab2),
           .a1b0_1sc(din_32_ab0_1sc), .a1b1_1sc(din_32_ab1_1sc), .a1b2_1sc(din_32_ab2_1sc),
           .msk_a1b0(din_32_msk_ab0), .msk_a1b1(din_32_msk_ab1), .msk_a1b2(din_32_msk_ab2),
           .msk_a1b0_1sc(din_32_msk_ab0_1sc), .msk_a1b1_1sc(din_32_msk_ab1_1sc), .msk_a1b2_1sc(din_32_msk_ab2_1sc),

           .a2b0(din_34_ab0), .a2b1(din_34_ab1),
           .a2b0_1sc(din_34_ab0_1sc), .a2b1_1sc(din_34_ab1_1sc),
           .msk_a2b0(din_34_msk_ab0), .msk_a2b1(din_34_msk_ab1),
           .msk_a2b0_1sc(din_34_msk_ab0_1sc), .msk_a2b1_1sc(din_34_msk_ab1_1sc),
           
           .a3b0(din_36_ab0),
           .a3b0_1sc(din_36_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12)
) addr_2_31_calc (
           .clk(clk), .sign(din_signs_reg[31]), 
           .p(addr_2_31),
           .a0b0(din_31_ab0), .a0b1(din_31_ab1), .a0b2(din_31_ab2), .a0b3(din_31_ab3),
           .a0b0_1sc(din_31_ab0_1sc), .a0b1_1sc(din_31_ab1_1sc), .a0b2_1sc(din_31_ab2_1sc), .a0b3_1sc(din_31_ab3_1sc),
           .msk_a0b0(din_31_msk_ab0), .msk_a0b1(din_31_msk_ab1), .msk_a0b2(din_31_msk_ab2), .msk_a0b3(din_31_msk_ab3),
           .msk_a0b0_1sc(din_31_msk_ab0_1sc), .msk_a0b1_1sc(din_31_msk_ab1_1sc), .msk_a0b2_1sc(din_31_msk_ab2_1sc), .msk_a0b3_1sc(din_31_msk_ab3_1sc),

           .a1b0(din_33_ab0), .a1b1(din_33_ab1), .a1b2(din_33_ab2),
           .a1b0_1sc(din_33_ab0_1sc), .a1b1_1sc(din_33_ab1_1sc), .a1b2_1sc(din_33_ab2_1sc),
           .msk_a1b0(din_33_msk_ab0), .msk_a1b1(din_33_msk_ab1), .msk_a1b2(din_33_msk_ab2),
           .msk_a1b0_1sc(din_33_msk_ab0_1sc), .msk_a1b1_1sc(din_33_msk_ab1_1sc), .msk_a1b2_1sc(din_33_msk_ab2_1sc),

           .a2b0(din_35_ab0), .a2b1(din_35_ab1),
           .a2b0_1sc(din_35_ab0_1sc), .a2b1_1sc(din_35_ab1_1sc),
           .msk_a2b0(din_35_msk_ab0), .msk_a2b1(din_35_msk_ab1),
           .msk_a2b0_1sc(din_35_msk_ab0_1sc), .msk_a2b1_1sc(din_35_msk_ab1_1sc),
           
           .a3b0(din_37_ab0),
           .a3b0_1sc(din_37_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_0_calc (
           .clk(clk), .sign(din_signs_reg[0]), 
           .p(addr_3_0),
           .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
           .a0b0_1sc(din_0_ab0_1sc), .a0b1_1sc(din_0_ab1_1sc), .a0b2_1sc(din_0_ab2_1sc), .a0b3_1sc(din_0_ab3_1sc),
           .msk_a0b0(din_0_msk_ab0), .msk_a0b1(din_0_msk_ab1), .msk_a0b2(din_0_msk_ab2), .msk_a0b3(din_0_msk_ab3),
           .msk_a0b0_1sc(din_0_msk_ab0_1sc), .msk_a0b1_1sc(din_0_msk_ab1_1sc), .msk_a0b2_1sc(din_0_msk_ab2_1sc), .msk_a0b3_1sc(din_0_msk_ab3_1sc),

           .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2),
           .a1b0_1sc(din_2_ab0_1sc), .a1b1_1sc(din_2_ab1_1sc), .a1b2_1sc(din_2_ab2_1sc),
           .msk_a1b0(din_2_msk_ab0), .msk_a1b1(din_2_msk_ab1), .msk_a1b2(din_2_msk_ab2),
           .msk_a1b0_1sc(din_2_msk_ab0_1sc), .msk_a1b1_1sc(din_2_msk_ab1_1sc), .msk_a1b2_1sc(din_2_msk_ab2_1sc),

           .a2b0(din_4_ab0), .a2b1(din_4_ab1),
           .a2b0_1sc(din_4_ab0_1sc), .a2b1_1sc(din_4_ab1_1sc),
           .msk_a2b0(din_4_msk_ab0), .msk_a2b1(din_4_msk_ab1),
           .msk_a2b0_1sc(din_4_msk_ab0_1sc), .msk_a2b1_1sc(din_4_msk_ab1_1sc),
           
           .a3b0(din_6_ab0),
           .a3b0_1sc(din_6_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_1_calc (
           .clk(clk), .sign(din_signs_reg[1]), 
           .p(addr_3_1),
           .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
           .a0b0_1sc(din_1_ab0_1sc), .a0b1_1sc(din_1_ab1_1sc), .a0b2_1sc(din_1_ab2_1sc), .a0b3_1sc(din_1_ab3_1sc),
           .msk_a0b0(din_1_msk_ab0), .msk_a0b1(din_1_msk_ab1), .msk_a0b2(din_1_msk_ab2), .msk_a0b3(din_1_msk_ab3),
           .msk_a0b0_1sc(din_1_msk_ab0_1sc), .msk_a0b1_1sc(din_1_msk_ab1_1sc), .msk_a0b2_1sc(din_1_msk_ab2_1sc), .msk_a0b3_1sc(din_1_msk_ab3_1sc),

           .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2),
           .a1b0_1sc(din_3_ab0_1sc), .a1b1_1sc(din_3_ab1_1sc), .a1b2_1sc(din_3_ab2_1sc),
           .msk_a1b0(din_3_msk_ab0), .msk_a1b1(din_3_msk_ab1), .msk_a1b2(din_3_msk_ab2),
           .msk_a1b0_1sc(din_3_msk_ab0_1sc), .msk_a1b1_1sc(din_3_msk_ab1_1sc), .msk_a1b2_1sc(din_3_msk_ab2_1sc),

           .a2b0(din_5_ab0), .a2b1(din_5_ab1),
           .a2b0_1sc(din_5_ab0_1sc), .a2b1_1sc(din_5_ab1_1sc),
           .msk_a2b0(din_5_msk_ab0), .msk_a2b1(din_5_msk_ab1),
           .msk_a2b0_1sc(din_5_msk_ab0_1sc), .msk_a2b1_1sc(din_5_msk_ab1_1sc),
           
           .a3b0(din_7_ab0),
           .a3b0_1sc(din_7_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_2_calc (
           .clk(clk), .sign(din_signs_reg[2]), 
           .p(addr_3_2),
           .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
           .a0b0_1sc(din_2_ab0_1sc), .a0b1_1sc(din_2_ab1_1sc), .a0b2_1sc(din_2_ab2_1sc), .a0b3_1sc(din_2_ab3_1sc),
           .msk_a0b0(din_2_msk_ab0), .msk_a0b1(din_2_msk_ab1), .msk_a0b2(din_2_msk_ab2), .msk_a0b3(din_2_msk_ab3),
           .msk_a0b0_1sc(din_2_msk_ab0_1sc), .msk_a0b1_1sc(din_2_msk_ab1_1sc), .msk_a0b2_1sc(din_2_msk_ab2_1sc), .msk_a0b3_1sc(din_2_msk_ab3_1sc),

           .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2),
           .a1b0_1sc(din_4_ab0_1sc), .a1b1_1sc(din_4_ab1_1sc), .a1b2_1sc(din_4_ab2_1sc),
           .msk_a1b0(din_4_msk_ab0), .msk_a1b1(din_4_msk_ab1), .msk_a1b2(din_4_msk_ab2),
           .msk_a1b0_1sc(din_4_msk_ab0_1sc), .msk_a1b1_1sc(din_4_msk_ab1_1sc), .msk_a1b2_1sc(din_4_msk_ab2_1sc),

           .a2b0(din_6_ab0), .a2b1(din_6_ab1),
           .a2b0_1sc(din_6_ab0_1sc), .a2b1_1sc(din_6_ab1_1sc),
           .msk_a2b0(din_6_msk_ab0), .msk_a2b1(din_6_msk_ab1),
           .msk_a2b0_1sc(din_6_msk_ab0_1sc), .msk_a2b1_1sc(din_6_msk_ab1_1sc),
           
           .a3b0(din_8_ab0),
           .a3b0_1sc(din_8_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_3_calc (
           .clk(clk), .sign(din_signs_reg[3]), 
           .p(addr_3_3),
           .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
           .a0b0_1sc(din_3_ab0_1sc), .a0b1_1sc(din_3_ab1_1sc), .a0b2_1sc(din_3_ab2_1sc), .a0b3_1sc(din_3_ab3_1sc),
           .msk_a0b0(din_3_msk_ab0), .msk_a0b1(din_3_msk_ab1), .msk_a0b2(din_3_msk_ab2), .msk_a0b3(din_3_msk_ab3),
           .msk_a0b0_1sc(din_3_msk_ab0_1sc), .msk_a0b1_1sc(din_3_msk_ab1_1sc), .msk_a0b2_1sc(din_3_msk_ab2_1sc), .msk_a0b3_1sc(din_3_msk_ab3_1sc),

           .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2),
           .a1b0_1sc(din_5_ab0_1sc), .a1b1_1sc(din_5_ab1_1sc), .a1b2_1sc(din_5_ab2_1sc),
           .msk_a1b0(din_5_msk_ab0), .msk_a1b1(din_5_msk_ab1), .msk_a1b2(din_5_msk_ab2),
           .msk_a1b0_1sc(din_5_msk_ab0_1sc), .msk_a1b1_1sc(din_5_msk_ab1_1sc), .msk_a1b2_1sc(din_5_msk_ab2_1sc),

           .a2b0(din_7_ab0), .a2b1(din_7_ab1),
           .a2b0_1sc(din_7_ab0_1sc), .a2b1_1sc(din_7_ab1_1sc),
           .msk_a2b0(din_7_msk_ab0), .msk_a2b1(din_7_msk_ab1),
           .msk_a2b0_1sc(din_7_msk_ab0_1sc), .msk_a2b1_1sc(din_7_msk_ab1_1sc),
           
           .a3b0(din_9_ab0),
           .a3b0_1sc(din_9_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_4_calc (
           .clk(clk), .sign(din_signs_reg[4]), 
           .p(addr_3_4),
           .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
           .a0b0_1sc(din_4_ab0_1sc), .a0b1_1sc(din_4_ab1_1sc), .a0b2_1sc(din_4_ab2_1sc), .a0b3_1sc(din_4_ab3_1sc),
           .msk_a0b0(din_4_msk_ab0), .msk_a0b1(din_4_msk_ab1), .msk_a0b2(din_4_msk_ab2), .msk_a0b3(din_4_msk_ab3),
           .msk_a0b0_1sc(din_4_msk_ab0_1sc), .msk_a0b1_1sc(din_4_msk_ab1_1sc), .msk_a0b2_1sc(din_4_msk_ab2_1sc), .msk_a0b3_1sc(din_4_msk_ab3_1sc),

           .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2),
           .a1b0_1sc(din_6_ab0_1sc), .a1b1_1sc(din_6_ab1_1sc), .a1b2_1sc(din_6_ab2_1sc),
           .msk_a1b0(din_6_msk_ab0), .msk_a1b1(din_6_msk_ab1), .msk_a1b2(din_6_msk_ab2),
           .msk_a1b0_1sc(din_6_msk_ab0_1sc), .msk_a1b1_1sc(din_6_msk_ab1_1sc), .msk_a1b2_1sc(din_6_msk_ab2_1sc),

           .a2b0(din_8_ab0), .a2b1(din_8_ab1),
           .a2b0_1sc(din_8_ab0_1sc), .a2b1_1sc(din_8_ab1_1sc),
           .msk_a2b0(din_8_msk_ab0), .msk_a2b1(din_8_msk_ab1),
           .msk_a2b0_1sc(din_8_msk_ab0_1sc), .msk_a2b1_1sc(din_8_msk_ab1_1sc),
           
           .a3b0(din_10_ab0),
           .a3b0_1sc(din_10_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_5_calc (
           .clk(clk), .sign(din_signs_reg[5]), 
           .p(addr_3_5),
           .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
           .a0b0_1sc(din_5_ab0_1sc), .a0b1_1sc(din_5_ab1_1sc), .a0b2_1sc(din_5_ab2_1sc), .a0b3_1sc(din_5_ab3_1sc),
           .msk_a0b0(din_5_msk_ab0), .msk_a0b1(din_5_msk_ab1), .msk_a0b2(din_5_msk_ab2), .msk_a0b3(din_5_msk_ab3),
           .msk_a0b0_1sc(din_5_msk_ab0_1sc), .msk_a0b1_1sc(din_5_msk_ab1_1sc), .msk_a0b2_1sc(din_5_msk_ab2_1sc), .msk_a0b3_1sc(din_5_msk_ab3_1sc),

           .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2),
           .a1b0_1sc(din_7_ab0_1sc), .a1b1_1sc(din_7_ab1_1sc), .a1b2_1sc(din_7_ab2_1sc),
           .msk_a1b0(din_7_msk_ab0), .msk_a1b1(din_7_msk_ab1), .msk_a1b2(din_7_msk_ab2),
           .msk_a1b0_1sc(din_7_msk_ab0_1sc), .msk_a1b1_1sc(din_7_msk_ab1_1sc), .msk_a1b2_1sc(din_7_msk_ab2_1sc),

           .a2b0(din_9_ab0), .a2b1(din_9_ab1),
           .a2b0_1sc(din_9_ab0_1sc), .a2b1_1sc(din_9_ab1_1sc),
           .msk_a2b0(din_9_msk_ab0), .msk_a2b1(din_9_msk_ab1),
           .msk_a2b0_1sc(din_9_msk_ab0_1sc), .msk_a2b1_1sc(din_9_msk_ab1_1sc),
           
           .a3b0(din_11_ab0),
           .a3b0_1sc(din_11_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_6_calc (
           .clk(clk), .sign(din_signs_reg[6]), 
           .p(addr_3_6),
           .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
           .a0b0_1sc(din_6_ab0_1sc), .a0b1_1sc(din_6_ab1_1sc), .a0b2_1sc(din_6_ab2_1sc), .a0b3_1sc(din_6_ab3_1sc),
           .msk_a0b0(din_6_msk_ab0), .msk_a0b1(din_6_msk_ab1), .msk_a0b2(din_6_msk_ab2), .msk_a0b3(din_6_msk_ab3),
           .msk_a0b0_1sc(din_6_msk_ab0_1sc), .msk_a0b1_1sc(din_6_msk_ab1_1sc), .msk_a0b2_1sc(din_6_msk_ab2_1sc), .msk_a0b3_1sc(din_6_msk_ab3_1sc),

           .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2),
           .a1b0_1sc(din_8_ab0_1sc), .a1b1_1sc(din_8_ab1_1sc), .a1b2_1sc(din_8_ab2_1sc),
           .msk_a1b0(din_8_msk_ab0), .msk_a1b1(din_8_msk_ab1), .msk_a1b2(din_8_msk_ab2),
           .msk_a1b0_1sc(din_8_msk_ab0_1sc), .msk_a1b1_1sc(din_8_msk_ab1_1sc), .msk_a1b2_1sc(din_8_msk_ab2_1sc),

           .a2b0(din_10_ab0), .a2b1(din_10_ab1),
           .a2b0_1sc(din_10_ab0_1sc), .a2b1_1sc(din_10_ab1_1sc),
           .msk_a2b0(din_10_msk_ab0), .msk_a2b1(din_10_msk_ab1),
           .msk_a2b0_1sc(din_10_msk_ab0_1sc), .msk_a2b1_1sc(din_10_msk_ab1_1sc),
           
           .a3b0(din_12_ab0),
           .a3b0_1sc(din_12_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_7_calc (
           .clk(clk), .sign(din_signs_reg[7]), 
           .p(addr_3_7),
           .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
           .a0b0_1sc(din_7_ab0_1sc), .a0b1_1sc(din_7_ab1_1sc), .a0b2_1sc(din_7_ab2_1sc), .a0b3_1sc(din_7_ab3_1sc),
           .msk_a0b0(din_7_msk_ab0), .msk_a0b1(din_7_msk_ab1), .msk_a0b2(din_7_msk_ab2), .msk_a0b3(din_7_msk_ab3),
           .msk_a0b0_1sc(din_7_msk_ab0_1sc), .msk_a0b1_1sc(din_7_msk_ab1_1sc), .msk_a0b2_1sc(din_7_msk_ab2_1sc), .msk_a0b3_1sc(din_7_msk_ab3_1sc),

           .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2),
           .a1b0_1sc(din_9_ab0_1sc), .a1b1_1sc(din_9_ab1_1sc), .a1b2_1sc(din_9_ab2_1sc),
           .msk_a1b0(din_9_msk_ab0), .msk_a1b1(din_9_msk_ab1), .msk_a1b2(din_9_msk_ab2),
           .msk_a1b0_1sc(din_9_msk_ab0_1sc), .msk_a1b1_1sc(din_9_msk_ab1_1sc), .msk_a1b2_1sc(din_9_msk_ab2_1sc),

           .a2b0(din_11_ab0), .a2b1(din_11_ab1),
           .a2b0_1sc(din_11_ab0_1sc), .a2b1_1sc(din_11_ab1_1sc),
           .msk_a2b0(din_11_msk_ab0), .msk_a2b1(din_11_msk_ab1),
           .msk_a2b0_1sc(din_11_msk_ab0_1sc), .msk_a2b1_1sc(din_11_msk_ab1_1sc),
           
           .a3b0(din_13_ab0),
           .a3b0_1sc(din_13_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_8_calc (
           .clk(clk), .sign(din_signs_reg[8]), 
           .p(addr_3_8),
           .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
           .a0b0_1sc(din_8_ab0_1sc), .a0b1_1sc(din_8_ab1_1sc), .a0b2_1sc(din_8_ab2_1sc), .a0b3_1sc(din_8_ab3_1sc),
           .msk_a0b0(din_8_msk_ab0), .msk_a0b1(din_8_msk_ab1), .msk_a0b2(din_8_msk_ab2), .msk_a0b3(din_8_msk_ab3),
           .msk_a0b0_1sc(din_8_msk_ab0_1sc), .msk_a0b1_1sc(din_8_msk_ab1_1sc), .msk_a0b2_1sc(din_8_msk_ab2_1sc), .msk_a0b3_1sc(din_8_msk_ab3_1sc),

           .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2),
           .a1b0_1sc(din_10_ab0_1sc), .a1b1_1sc(din_10_ab1_1sc), .a1b2_1sc(din_10_ab2_1sc),
           .msk_a1b0(din_10_msk_ab0), .msk_a1b1(din_10_msk_ab1), .msk_a1b2(din_10_msk_ab2),
           .msk_a1b0_1sc(din_10_msk_ab0_1sc), .msk_a1b1_1sc(din_10_msk_ab1_1sc), .msk_a1b2_1sc(din_10_msk_ab2_1sc),

           .a2b0(din_12_ab0), .a2b1(din_12_ab1),
           .a2b0_1sc(din_12_ab0_1sc), .a2b1_1sc(din_12_ab1_1sc),
           .msk_a2b0(din_12_msk_ab0), .msk_a2b1(din_12_msk_ab1),
           .msk_a2b0_1sc(din_12_msk_ab0_1sc), .msk_a2b1_1sc(din_12_msk_ab1_1sc),
           
           .a3b0(din_14_ab0),
           .a3b0_1sc(din_14_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_9_calc (
           .clk(clk), .sign(din_signs_reg[9]), 
           .p(addr_3_9),
           .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
           .a0b0_1sc(din_9_ab0_1sc), .a0b1_1sc(din_9_ab1_1sc), .a0b2_1sc(din_9_ab2_1sc), .a0b3_1sc(din_9_ab3_1sc),
           .msk_a0b0(din_9_msk_ab0), .msk_a0b1(din_9_msk_ab1), .msk_a0b2(din_9_msk_ab2), .msk_a0b3(din_9_msk_ab3),
           .msk_a0b0_1sc(din_9_msk_ab0_1sc), .msk_a0b1_1sc(din_9_msk_ab1_1sc), .msk_a0b2_1sc(din_9_msk_ab2_1sc), .msk_a0b3_1sc(din_9_msk_ab3_1sc),

           .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2),
           .a1b0_1sc(din_11_ab0_1sc), .a1b1_1sc(din_11_ab1_1sc), .a1b2_1sc(din_11_ab2_1sc),
           .msk_a1b0(din_11_msk_ab0), .msk_a1b1(din_11_msk_ab1), .msk_a1b2(din_11_msk_ab2),
           .msk_a1b0_1sc(din_11_msk_ab0_1sc), .msk_a1b1_1sc(din_11_msk_ab1_1sc), .msk_a1b2_1sc(din_11_msk_ab2_1sc),

           .a2b0(din_13_ab0), .a2b1(din_13_ab1),
           .a2b0_1sc(din_13_ab0_1sc), .a2b1_1sc(din_13_ab1_1sc),
           .msk_a2b0(din_13_msk_ab0), .msk_a2b1(din_13_msk_ab1),
           .msk_a2b0_1sc(din_13_msk_ab0_1sc), .msk_a2b1_1sc(din_13_msk_ab1_1sc),
           
           .a3b0(din_15_ab0),
           .a3b0_1sc(din_15_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_10_calc (
           .clk(clk), .sign(din_signs_reg[10]), 
           .p(addr_3_10),
           .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
           .a0b0_1sc(din_10_ab0_1sc), .a0b1_1sc(din_10_ab1_1sc), .a0b2_1sc(din_10_ab2_1sc), .a0b3_1sc(din_10_ab3_1sc),
           .msk_a0b0(din_10_msk_ab0), .msk_a0b1(din_10_msk_ab1), .msk_a0b2(din_10_msk_ab2), .msk_a0b3(din_10_msk_ab3),
           .msk_a0b0_1sc(din_10_msk_ab0_1sc), .msk_a0b1_1sc(din_10_msk_ab1_1sc), .msk_a0b2_1sc(din_10_msk_ab2_1sc), .msk_a0b3_1sc(din_10_msk_ab3_1sc),

           .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2),
           .a1b0_1sc(din_12_ab0_1sc), .a1b1_1sc(din_12_ab1_1sc), .a1b2_1sc(din_12_ab2_1sc),
           .msk_a1b0(din_12_msk_ab0), .msk_a1b1(din_12_msk_ab1), .msk_a1b2(din_12_msk_ab2),
           .msk_a1b0_1sc(din_12_msk_ab0_1sc), .msk_a1b1_1sc(din_12_msk_ab1_1sc), .msk_a1b2_1sc(din_12_msk_ab2_1sc),

           .a2b0(din_14_ab0), .a2b1(din_14_ab1),
           .a2b0_1sc(din_14_ab0_1sc), .a2b1_1sc(din_14_ab1_1sc),
           .msk_a2b0(din_14_msk_ab0), .msk_a2b1(din_14_msk_ab1),
           .msk_a2b0_1sc(din_14_msk_ab0_1sc), .msk_a2b1_1sc(din_14_msk_ab1_1sc),
           
           .a3b0(din_16_ab0),
           .a3b0_1sc(din_16_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_11_calc (
           .clk(clk), .sign(din_signs_reg[11]), 
           .p(addr_3_11),
           .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
           .a0b0_1sc(din_11_ab0_1sc), .a0b1_1sc(din_11_ab1_1sc), .a0b2_1sc(din_11_ab2_1sc), .a0b3_1sc(din_11_ab3_1sc),
           .msk_a0b0(din_11_msk_ab0), .msk_a0b1(din_11_msk_ab1), .msk_a0b2(din_11_msk_ab2), .msk_a0b3(din_11_msk_ab3),
           .msk_a0b0_1sc(din_11_msk_ab0_1sc), .msk_a0b1_1sc(din_11_msk_ab1_1sc), .msk_a0b2_1sc(din_11_msk_ab2_1sc), .msk_a0b3_1sc(din_11_msk_ab3_1sc),

           .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2),
           .a1b0_1sc(din_13_ab0_1sc), .a1b1_1sc(din_13_ab1_1sc), .a1b2_1sc(din_13_ab2_1sc),
           .msk_a1b0(din_13_msk_ab0), .msk_a1b1(din_13_msk_ab1), .msk_a1b2(din_13_msk_ab2),
           .msk_a1b0_1sc(din_13_msk_ab0_1sc), .msk_a1b1_1sc(din_13_msk_ab1_1sc), .msk_a1b2_1sc(din_13_msk_ab2_1sc),

           .a2b0(din_15_ab0), .a2b1(din_15_ab1),
           .a2b0_1sc(din_15_ab0_1sc), .a2b1_1sc(din_15_ab1_1sc),
           .msk_a2b0(din_15_msk_ab0), .msk_a2b1(din_15_msk_ab1),
           .msk_a2b0_1sc(din_15_msk_ab0_1sc), .msk_a2b1_1sc(din_15_msk_ab1_1sc),
           
           .a3b0(din_17_ab0),
           .a3b0_1sc(din_17_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_12_calc (
           .clk(clk), .sign(din_signs_reg[12]), 
           .p(addr_3_12),
           .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
           .a0b0_1sc(din_12_ab0_1sc), .a0b1_1sc(din_12_ab1_1sc), .a0b2_1sc(din_12_ab2_1sc), .a0b3_1sc(din_12_ab3_1sc),
           .msk_a0b0(din_12_msk_ab0), .msk_a0b1(din_12_msk_ab1), .msk_a0b2(din_12_msk_ab2), .msk_a0b3(din_12_msk_ab3),
           .msk_a0b0_1sc(din_12_msk_ab0_1sc), .msk_a0b1_1sc(din_12_msk_ab1_1sc), .msk_a0b2_1sc(din_12_msk_ab2_1sc), .msk_a0b3_1sc(din_12_msk_ab3_1sc),

           .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2),
           .a1b0_1sc(din_14_ab0_1sc), .a1b1_1sc(din_14_ab1_1sc), .a1b2_1sc(din_14_ab2_1sc),
           .msk_a1b0(din_14_msk_ab0), .msk_a1b1(din_14_msk_ab1), .msk_a1b2(din_14_msk_ab2),
           .msk_a1b0_1sc(din_14_msk_ab0_1sc), .msk_a1b1_1sc(din_14_msk_ab1_1sc), .msk_a1b2_1sc(din_14_msk_ab2_1sc),

           .a2b0(din_16_ab0), .a2b1(din_16_ab1),
           .a2b0_1sc(din_16_ab0_1sc), .a2b1_1sc(din_16_ab1_1sc),
           .msk_a2b0(din_16_msk_ab0), .msk_a2b1(din_16_msk_ab1),
           .msk_a2b0_1sc(din_16_msk_ab0_1sc), .msk_a2b1_1sc(din_16_msk_ab1_1sc),
           
           .a3b0(din_18_ab0),
           .a3b0_1sc(din_18_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_13_calc (
           .clk(clk), .sign(din_signs_reg[13]), 
           .p(addr_3_13),
           .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
           .a0b0_1sc(din_13_ab0_1sc), .a0b1_1sc(din_13_ab1_1sc), .a0b2_1sc(din_13_ab2_1sc), .a0b3_1sc(din_13_ab3_1sc),
           .msk_a0b0(din_13_msk_ab0), .msk_a0b1(din_13_msk_ab1), .msk_a0b2(din_13_msk_ab2), .msk_a0b3(din_13_msk_ab3),
           .msk_a0b0_1sc(din_13_msk_ab0_1sc), .msk_a0b1_1sc(din_13_msk_ab1_1sc), .msk_a0b2_1sc(din_13_msk_ab2_1sc), .msk_a0b3_1sc(din_13_msk_ab3_1sc),

           .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2),
           .a1b0_1sc(din_15_ab0_1sc), .a1b1_1sc(din_15_ab1_1sc), .a1b2_1sc(din_15_ab2_1sc),
           .msk_a1b0(din_15_msk_ab0), .msk_a1b1(din_15_msk_ab1), .msk_a1b2(din_15_msk_ab2),
           .msk_a1b0_1sc(din_15_msk_ab0_1sc), .msk_a1b1_1sc(din_15_msk_ab1_1sc), .msk_a1b2_1sc(din_15_msk_ab2_1sc),

           .a2b0(din_17_ab0), .a2b1(din_17_ab1),
           .a2b0_1sc(din_17_ab0_1sc), .a2b1_1sc(din_17_ab1_1sc),
           .msk_a2b0(din_17_msk_ab0), .msk_a2b1(din_17_msk_ab1),
           .msk_a2b0_1sc(din_17_msk_ab0_1sc), .msk_a2b1_1sc(din_17_msk_ab1_1sc),
           
           .a3b0(din_19_ab0),
           .a3b0_1sc(din_19_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_14_calc (
           .clk(clk), .sign(din_signs_reg[14]), 
           .p(addr_3_14),
           .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
           .a0b0_1sc(din_14_ab0_1sc), .a0b1_1sc(din_14_ab1_1sc), .a0b2_1sc(din_14_ab2_1sc), .a0b3_1sc(din_14_ab3_1sc),
           .msk_a0b0(din_14_msk_ab0), .msk_a0b1(din_14_msk_ab1), .msk_a0b2(din_14_msk_ab2), .msk_a0b3(din_14_msk_ab3),
           .msk_a0b0_1sc(din_14_msk_ab0_1sc), .msk_a0b1_1sc(din_14_msk_ab1_1sc), .msk_a0b2_1sc(din_14_msk_ab2_1sc), .msk_a0b3_1sc(din_14_msk_ab3_1sc),

           .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2),
           .a1b0_1sc(din_16_ab0_1sc), .a1b1_1sc(din_16_ab1_1sc), .a1b2_1sc(din_16_ab2_1sc),
           .msk_a1b0(din_16_msk_ab0), .msk_a1b1(din_16_msk_ab1), .msk_a1b2(din_16_msk_ab2),
           .msk_a1b0_1sc(din_16_msk_ab0_1sc), .msk_a1b1_1sc(din_16_msk_ab1_1sc), .msk_a1b2_1sc(din_16_msk_ab2_1sc),

           .a2b0(din_18_ab0), .a2b1(din_18_ab1),
           .a2b0_1sc(din_18_ab0_1sc), .a2b1_1sc(din_18_ab1_1sc),
           .msk_a2b0(din_18_msk_ab0), .msk_a2b1(din_18_msk_ab1),
           .msk_a2b0_1sc(din_18_msk_ab0_1sc), .msk_a2b1_1sc(din_18_msk_ab1_1sc),
           
           .a3b0(din_20_ab0),
           .a3b0_1sc(din_20_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_15_calc (
           .clk(clk), .sign(din_signs_reg[15]), 
           .p(addr_3_15),
           .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
           .a0b0_1sc(din_15_ab0_1sc), .a0b1_1sc(din_15_ab1_1sc), .a0b2_1sc(din_15_ab2_1sc), .a0b3_1sc(din_15_ab3_1sc),
           .msk_a0b0(din_15_msk_ab0), .msk_a0b1(din_15_msk_ab1), .msk_a0b2(din_15_msk_ab2), .msk_a0b3(din_15_msk_ab3),
           .msk_a0b0_1sc(din_15_msk_ab0_1sc), .msk_a0b1_1sc(din_15_msk_ab1_1sc), .msk_a0b2_1sc(din_15_msk_ab2_1sc), .msk_a0b3_1sc(din_15_msk_ab3_1sc),

           .a1b0(din_17_ab0), .a1b1(din_17_ab1), .a1b2(din_17_ab2),
           .a1b0_1sc(din_17_ab0_1sc), .a1b1_1sc(din_17_ab1_1sc), .a1b2_1sc(din_17_ab2_1sc),
           .msk_a1b0(din_17_msk_ab0), .msk_a1b1(din_17_msk_ab1), .msk_a1b2(din_17_msk_ab2),
           .msk_a1b0_1sc(din_17_msk_ab0_1sc), .msk_a1b1_1sc(din_17_msk_ab1_1sc), .msk_a1b2_1sc(din_17_msk_ab2_1sc),

           .a2b0(din_19_ab0), .a2b1(din_19_ab1),
           .a2b0_1sc(din_19_ab0_1sc), .a2b1_1sc(din_19_ab1_1sc),
           .msk_a2b0(din_19_msk_ab0), .msk_a2b1(din_19_msk_ab1),
           .msk_a2b0_1sc(din_19_msk_ab0_1sc), .msk_a2b1_1sc(din_19_msk_ab1_1sc),
           
           .a3b0(din_21_ab0),
           .a3b0_1sc(din_21_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_16_calc (
           .clk(clk), .sign(din_signs_reg[16]), 
           .p(addr_3_16),
           .a0b0(din_16_ab0), .a0b1(din_16_ab1), .a0b2(din_16_ab2), .a0b3(din_16_ab3),
           .a0b0_1sc(din_16_ab0_1sc), .a0b1_1sc(din_16_ab1_1sc), .a0b2_1sc(din_16_ab2_1sc), .a0b3_1sc(din_16_ab3_1sc),
           .msk_a0b0(din_16_msk_ab0), .msk_a0b1(din_16_msk_ab1), .msk_a0b2(din_16_msk_ab2), .msk_a0b3(din_16_msk_ab3),
           .msk_a0b0_1sc(din_16_msk_ab0_1sc), .msk_a0b1_1sc(din_16_msk_ab1_1sc), .msk_a0b2_1sc(din_16_msk_ab2_1sc), .msk_a0b3_1sc(din_16_msk_ab3_1sc),

           .a1b0(din_18_ab0), .a1b1(din_18_ab1), .a1b2(din_18_ab2),
           .a1b0_1sc(din_18_ab0_1sc), .a1b1_1sc(din_18_ab1_1sc), .a1b2_1sc(din_18_ab2_1sc),
           .msk_a1b0(din_18_msk_ab0), .msk_a1b1(din_18_msk_ab1), .msk_a1b2(din_18_msk_ab2),
           .msk_a1b0_1sc(din_18_msk_ab0_1sc), .msk_a1b1_1sc(din_18_msk_ab1_1sc), .msk_a1b2_1sc(din_18_msk_ab2_1sc),

           .a2b0(din_20_ab0), .a2b1(din_20_ab1),
           .a2b0_1sc(din_20_ab0_1sc), .a2b1_1sc(din_20_ab1_1sc),
           .msk_a2b0(din_20_msk_ab0), .msk_a2b1(din_20_msk_ab1),
           .msk_a2b0_1sc(din_20_msk_ab0_1sc), .msk_a2b1_1sc(din_20_msk_ab1_1sc),
           
           .a3b0(din_22_ab0),
           .a3b0_1sc(din_22_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_17_calc (
           .clk(clk), .sign(din_signs_reg[17]), 
           .p(addr_3_17),
           .a0b0(din_17_ab0), .a0b1(din_17_ab1), .a0b2(din_17_ab2), .a0b3(din_17_ab3),
           .a0b0_1sc(din_17_ab0_1sc), .a0b1_1sc(din_17_ab1_1sc), .a0b2_1sc(din_17_ab2_1sc), .a0b3_1sc(din_17_ab3_1sc),
           .msk_a0b0(din_17_msk_ab0), .msk_a0b1(din_17_msk_ab1), .msk_a0b2(din_17_msk_ab2), .msk_a0b3(din_17_msk_ab3),
           .msk_a0b0_1sc(din_17_msk_ab0_1sc), .msk_a0b1_1sc(din_17_msk_ab1_1sc), .msk_a0b2_1sc(din_17_msk_ab2_1sc), .msk_a0b3_1sc(din_17_msk_ab3_1sc),

           .a1b0(din_19_ab0), .a1b1(din_19_ab1), .a1b2(din_19_ab2),
           .a1b0_1sc(din_19_ab0_1sc), .a1b1_1sc(din_19_ab1_1sc), .a1b2_1sc(din_19_ab2_1sc),
           .msk_a1b0(din_19_msk_ab0), .msk_a1b1(din_19_msk_ab1), .msk_a1b2(din_19_msk_ab2),
           .msk_a1b0_1sc(din_19_msk_ab0_1sc), .msk_a1b1_1sc(din_19_msk_ab1_1sc), .msk_a1b2_1sc(din_19_msk_ab2_1sc),

           .a2b0(din_21_ab0), .a2b1(din_21_ab1),
           .a2b0_1sc(din_21_ab0_1sc), .a2b1_1sc(din_21_ab1_1sc),
           .msk_a2b0(din_21_msk_ab0), .msk_a2b1(din_21_msk_ab1),
           .msk_a2b0_1sc(din_21_msk_ab0_1sc), .msk_a2b1_1sc(din_21_msk_ab1_1sc),
           
           .a3b0(din_23_ab0),
           .a3b0_1sc(din_23_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_18_calc (
           .clk(clk), .sign(din_signs_reg[18]), 
           .p(addr_3_18),
           .a0b0(din_18_ab0), .a0b1(din_18_ab1), .a0b2(din_18_ab2), .a0b3(din_18_ab3),
           .a0b0_1sc(din_18_ab0_1sc), .a0b1_1sc(din_18_ab1_1sc), .a0b2_1sc(din_18_ab2_1sc), .a0b3_1sc(din_18_ab3_1sc),
           .msk_a0b0(din_18_msk_ab0), .msk_a0b1(din_18_msk_ab1), .msk_a0b2(din_18_msk_ab2), .msk_a0b3(din_18_msk_ab3),
           .msk_a0b0_1sc(din_18_msk_ab0_1sc), .msk_a0b1_1sc(din_18_msk_ab1_1sc), .msk_a0b2_1sc(din_18_msk_ab2_1sc), .msk_a0b3_1sc(din_18_msk_ab3_1sc),

           .a1b0(din_20_ab0), .a1b1(din_20_ab1), .a1b2(din_20_ab2),
           .a1b0_1sc(din_20_ab0_1sc), .a1b1_1sc(din_20_ab1_1sc), .a1b2_1sc(din_20_ab2_1sc),
           .msk_a1b0(din_20_msk_ab0), .msk_a1b1(din_20_msk_ab1), .msk_a1b2(din_20_msk_ab2),
           .msk_a1b0_1sc(din_20_msk_ab0_1sc), .msk_a1b1_1sc(din_20_msk_ab1_1sc), .msk_a1b2_1sc(din_20_msk_ab2_1sc),

           .a2b0(din_22_ab0), .a2b1(din_22_ab1),
           .a2b0_1sc(din_22_ab0_1sc), .a2b1_1sc(din_22_ab1_1sc),
           .msk_a2b0(din_22_msk_ab0), .msk_a2b1(din_22_msk_ab1),
           .msk_a2b0_1sc(din_22_msk_ab0_1sc), .msk_a2b1_1sc(din_22_msk_ab1_1sc),
           
           .a3b0(din_24_ab0),
           .a3b0_1sc(din_24_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_19_calc (
           .clk(clk), .sign(din_signs_reg[19]), 
           .p(addr_3_19),
           .a0b0(din_19_ab0), .a0b1(din_19_ab1), .a0b2(din_19_ab2), .a0b3(din_19_ab3),
           .a0b0_1sc(din_19_ab0_1sc), .a0b1_1sc(din_19_ab1_1sc), .a0b2_1sc(din_19_ab2_1sc), .a0b3_1sc(din_19_ab3_1sc),
           .msk_a0b0(din_19_msk_ab0), .msk_a0b1(din_19_msk_ab1), .msk_a0b2(din_19_msk_ab2), .msk_a0b3(din_19_msk_ab3),
           .msk_a0b0_1sc(din_19_msk_ab0_1sc), .msk_a0b1_1sc(din_19_msk_ab1_1sc), .msk_a0b2_1sc(din_19_msk_ab2_1sc), .msk_a0b3_1sc(din_19_msk_ab3_1sc),

           .a1b0(din_21_ab0), .a1b1(din_21_ab1), .a1b2(din_21_ab2),
           .a1b0_1sc(din_21_ab0_1sc), .a1b1_1sc(din_21_ab1_1sc), .a1b2_1sc(din_21_ab2_1sc),
           .msk_a1b0(din_21_msk_ab0), .msk_a1b1(din_21_msk_ab1), .msk_a1b2(din_21_msk_ab2),
           .msk_a1b0_1sc(din_21_msk_ab0_1sc), .msk_a1b1_1sc(din_21_msk_ab1_1sc), .msk_a1b2_1sc(din_21_msk_ab2_1sc),

           .a2b0(din_23_ab0), .a2b1(din_23_ab1),
           .a2b0_1sc(din_23_ab0_1sc), .a2b1_1sc(din_23_ab1_1sc),
           .msk_a2b0(din_23_msk_ab0), .msk_a2b1(din_23_msk_ab1),
           .msk_a2b0_1sc(din_23_msk_ab0_1sc), .msk_a2b1_1sc(din_23_msk_ab1_1sc),
           
           .a3b0(din_25_ab0),
           .a3b0_1sc(din_25_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_20_calc (
           .clk(clk), .sign(din_signs_reg[20]), 
           .p(addr_3_20),
           .a0b0(din_20_ab0), .a0b1(din_20_ab1), .a0b2(din_20_ab2), .a0b3(din_20_ab3),
           .a0b0_1sc(din_20_ab0_1sc), .a0b1_1sc(din_20_ab1_1sc), .a0b2_1sc(din_20_ab2_1sc), .a0b3_1sc(din_20_ab3_1sc),
           .msk_a0b0(din_20_msk_ab0), .msk_a0b1(din_20_msk_ab1), .msk_a0b2(din_20_msk_ab2), .msk_a0b3(din_20_msk_ab3),
           .msk_a0b0_1sc(din_20_msk_ab0_1sc), .msk_a0b1_1sc(din_20_msk_ab1_1sc), .msk_a0b2_1sc(din_20_msk_ab2_1sc), .msk_a0b3_1sc(din_20_msk_ab3_1sc),

           .a1b0(din_22_ab0), .a1b1(din_22_ab1), .a1b2(din_22_ab2),
           .a1b0_1sc(din_22_ab0_1sc), .a1b1_1sc(din_22_ab1_1sc), .a1b2_1sc(din_22_ab2_1sc),
           .msk_a1b0(din_22_msk_ab0), .msk_a1b1(din_22_msk_ab1), .msk_a1b2(din_22_msk_ab2),
           .msk_a1b0_1sc(din_22_msk_ab0_1sc), .msk_a1b1_1sc(din_22_msk_ab1_1sc), .msk_a1b2_1sc(din_22_msk_ab2_1sc),

           .a2b0(din_24_ab0), .a2b1(din_24_ab1),
           .a2b0_1sc(din_24_ab0_1sc), .a2b1_1sc(din_24_ab1_1sc),
           .msk_a2b0(din_24_msk_ab0), .msk_a2b1(din_24_msk_ab1),
           .msk_a2b0_1sc(din_24_msk_ab0_1sc), .msk_a2b1_1sc(din_24_msk_ab1_1sc),
           
           .a3b0(din_26_ab0),
           .a3b0_1sc(din_26_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_21_calc (
           .clk(clk), .sign(din_signs_reg[21]), 
           .p(addr_3_21),
           .a0b0(din_21_ab0), .a0b1(din_21_ab1), .a0b2(din_21_ab2), .a0b3(din_21_ab3),
           .a0b0_1sc(din_21_ab0_1sc), .a0b1_1sc(din_21_ab1_1sc), .a0b2_1sc(din_21_ab2_1sc), .a0b3_1sc(din_21_ab3_1sc),
           .msk_a0b0(din_21_msk_ab0), .msk_a0b1(din_21_msk_ab1), .msk_a0b2(din_21_msk_ab2), .msk_a0b3(din_21_msk_ab3),
           .msk_a0b0_1sc(din_21_msk_ab0_1sc), .msk_a0b1_1sc(din_21_msk_ab1_1sc), .msk_a0b2_1sc(din_21_msk_ab2_1sc), .msk_a0b3_1sc(din_21_msk_ab3_1sc),

           .a1b0(din_23_ab0), .a1b1(din_23_ab1), .a1b2(din_23_ab2),
           .a1b0_1sc(din_23_ab0_1sc), .a1b1_1sc(din_23_ab1_1sc), .a1b2_1sc(din_23_ab2_1sc),
           .msk_a1b0(din_23_msk_ab0), .msk_a1b1(din_23_msk_ab1), .msk_a1b2(din_23_msk_ab2),
           .msk_a1b0_1sc(din_23_msk_ab0_1sc), .msk_a1b1_1sc(din_23_msk_ab1_1sc), .msk_a1b2_1sc(din_23_msk_ab2_1sc),

           .a2b0(din_25_ab0), .a2b1(din_25_ab1),
           .a2b0_1sc(din_25_ab0_1sc), .a2b1_1sc(din_25_ab1_1sc),
           .msk_a2b0(din_25_msk_ab0), .msk_a2b1(din_25_msk_ab1),
           .msk_a2b0_1sc(din_25_msk_ab0_1sc), .msk_a2b1_1sc(din_25_msk_ab1_1sc),
           
           .a3b0(din_27_ab0),
           .a3b0_1sc(din_27_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_22_calc (
           .clk(clk), .sign(din_signs_reg[22]), 
           .p(addr_3_22),
           .a0b0(din_22_ab0), .a0b1(din_22_ab1), .a0b2(din_22_ab2), .a0b3(din_22_ab3),
           .a0b0_1sc(din_22_ab0_1sc), .a0b1_1sc(din_22_ab1_1sc), .a0b2_1sc(din_22_ab2_1sc), .a0b3_1sc(din_22_ab3_1sc),
           .msk_a0b0(din_22_msk_ab0), .msk_a0b1(din_22_msk_ab1), .msk_a0b2(din_22_msk_ab2), .msk_a0b3(din_22_msk_ab3),
           .msk_a0b0_1sc(din_22_msk_ab0_1sc), .msk_a0b1_1sc(din_22_msk_ab1_1sc), .msk_a0b2_1sc(din_22_msk_ab2_1sc), .msk_a0b3_1sc(din_22_msk_ab3_1sc),

           .a1b0(din_24_ab0), .a1b1(din_24_ab1), .a1b2(din_24_ab2),
           .a1b0_1sc(din_24_ab0_1sc), .a1b1_1sc(din_24_ab1_1sc), .a1b2_1sc(din_24_ab2_1sc),
           .msk_a1b0(din_24_msk_ab0), .msk_a1b1(din_24_msk_ab1), .msk_a1b2(din_24_msk_ab2),
           .msk_a1b0_1sc(din_24_msk_ab0_1sc), .msk_a1b1_1sc(din_24_msk_ab1_1sc), .msk_a1b2_1sc(din_24_msk_ab2_1sc),

           .a2b0(din_26_ab0), .a2b1(din_26_ab1),
           .a2b0_1sc(din_26_ab0_1sc), .a2b1_1sc(din_26_ab1_1sc),
           .msk_a2b0(din_26_msk_ab0), .msk_a2b1(din_26_msk_ab1),
           .msk_a2b0_1sc(din_26_msk_ab0_1sc), .msk_a2b1_1sc(din_26_msk_ab1_1sc),
           
           .a3b0(din_28_ab0),
           .a3b0_1sc(din_28_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_23_calc (
           .clk(clk), .sign(din_signs_reg[23]), 
           .p(addr_3_23),
           .a0b0(din_23_ab0), .a0b1(din_23_ab1), .a0b2(din_23_ab2), .a0b3(din_23_ab3),
           .a0b0_1sc(din_23_ab0_1sc), .a0b1_1sc(din_23_ab1_1sc), .a0b2_1sc(din_23_ab2_1sc), .a0b3_1sc(din_23_ab3_1sc),
           .msk_a0b0(din_23_msk_ab0), .msk_a0b1(din_23_msk_ab1), .msk_a0b2(din_23_msk_ab2), .msk_a0b3(din_23_msk_ab3),
           .msk_a0b0_1sc(din_23_msk_ab0_1sc), .msk_a0b1_1sc(din_23_msk_ab1_1sc), .msk_a0b2_1sc(din_23_msk_ab2_1sc), .msk_a0b3_1sc(din_23_msk_ab3_1sc),

           .a1b0(din_25_ab0), .a1b1(din_25_ab1), .a1b2(din_25_ab2),
           .a1b0_1sc(din_25_ab0_1sc), .a1b1_1sc(din_25_ab1_1sc), .a1b2_1sc(din_25_ab2_1sc),
           .msk_a1b0(din_25_msk_ab0), .msk_a1b1(din_25_msk_ab1), .msk_a1b2(din_25_msk_ab2),
           .msk_a1b0_1sc(din_25_msk_ab0_1sc), .msk_a1b1_1sc(din_25_msk_ab1_1sc), .msk_a1b2_1sc(din_25_msk_ab2_1sc),

           .a2b0(din_27_ab0), .a2b1(din_27_ab1),
           .a2b0_1sc(din_27_ab0_1sc), .a2b1_1sc(din_27_ab1_1sc),
           .msk_a2b0(din_27_msk_ab0), .msk_a2b1(din_27_msk_ab1),
           .msk_a2b0_1sc(din_27_msk_ab0_1sc), .msk_a2b1_1sc(din_27_msk_ab1_1sc),
           
           .a3b0(din_29_ab0),
           .a3b0_1sc(din_29_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_24_calc (
           .clk(clk), .sign(din_signs_reg[24]), 
           .p(addr_3_24),
           .a0b0(din_24_ab0), .a0b1(din_24_ab1), .a0b2(din_24_ab2), .a0b3(din_24_ab3),
           .a0b0_1sc(din_24_ab0_1sc), .a0b1_1sc(din_24_ab1_1sc), .a0b2_1sc(din_24_ab2_1sc), .a0b3_1sc(din_24_ab3_1sc),
           .msk_a0b0(din_24_msk_ab0), .msk_a0b1(din_24_msk_ab1), .msk_a0b2(din_24_msk_ab2), .msk_a0b3(din_24_msk_ab3),
           .msk_a0b0_1sc(din_24_msk_ab0_1sc), .msk_a0b1_1sc(din_24_msk_ab1_1sc), .msk_a0b2_1sc(din_24_msk_ab2_1sc), .msk_a0b3_1sc(din_24_msk_ab3_1sc),

           .a1b0(din_26_ab0), .a1b1(din_26_ab1), .a1b2(din_26_ab2),
           .a1b0_1sc(din_26_ab0_1sc), .a1b1_1sc(din_26_ab1_1sc), .a1b2_1sc(din_26_ab2_1sc),
           .msk_a1b0(din_26_msk_ab0), .msk_a1b1(din_26_msk_ab1), .msk_a1b2(din_26_msk_ab2),
           .msk_a1b0_1sc(din_26_msk_ab0_1sc), .msk_a1b1_1sc(din_26_msk_ab1_1sc), .msk_a1b2_1sc(din_26_msk_ab2_1sc),

           .a2b0(din_28_ab0), .a2b1(din_28_ab1),
           .a2b0_1sc(din_28_ab0_1sc), .a2b1_1sc(din_28_ab1_1sc),
           .msk_a2b0(din_28_msk_ab0), .msk_a2b1(din_28_msk_ab1),
           .msk_a2b0_1sc(din_28_msk_ab0_1sc), .msk_a2b1_1sc(din_28_msk_ab1_1sc),
           
           .a3b0(din_30_ab0),
           .a3b0_1sc(din_30_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_25_calc (
           .clk(clk), .sign(din_signs_reg[25]), 
           .p(addr_3_25),
           .a0b0(din_25_ab0), .a0b1(din_25_ab1), .a0b2(din_25_ab2), .a0b3(din_25_ab3),
           .a0b0_1sc(din_25_ab0_1sc), .a0b1_1sc(din_25_ab1_1sc), .a0b2_1sc(din_25_ab2_1sc), .a0b3_1sc(din_25_ab3_1sc),
           .msk_a0b0(din_25_msk_ab0), .msk_a0b1(din_25_msk_ab1), .msk_a0b2(din_25_msk_ab2), .msk_a0b3(din_25_msk_ab3),
           .msk_a0b0_1sc(din_25_msk_ab0_1sc), .msk_a0b1_1sc(din_25_msk_ab1_1sc), .msk_a0b2_1sc(din_25_msk_ab2_1sc), .msk_a0b3_1sc(din_25_msk_ab3_1sc),

           .a1b0(din_27_ab0), .a1b1(din_27_ab1), .a1b2(din_27_ab2),
           .a1b0_1sc(din_27_ab0_1sc), .a1b1_1sc(din_27_ab1_1sc), .a1b2_1sc(din_27_ab2_1sc),
           .msk_a1b0(din_27_msk_ab0), .msk_a1b1(din_27_msk_ab1), .msk_a1b2(din_27_msk_ab2),
           .msk_a1b0_1sc(din_27_msk_ab0_1sc), .msk_a1b1_1sc(din_27_msk_ab1_1sc), .msk_a1b2_1sc(din_27_msk_ab2_1sc),

           .a2b0(din_29_ab0), .a2b1(din_29_ab1),
           .a2b0_1sc(din_29_ab0_1sc), .a2b1_1sc(din_29_ab1_1sc),
           .msk_a2b0(din_29_msk_ab0), .msk_a2b1(din_29_msk_ab1),
           .msk_a2b0_1sc(din_29_msk_ab0_1sc), .msk_a2b1_1sc(din_29_msk_ab1_1sc),
           
           .a3b0(din_31_ab0),
           .a3b0_1sc(din_31_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_26_calc (
           .clk(clk), .sign(din_signs_reg[26]), 
           .p(addr_3_26),
           .a0b0(din_26_ab0), .a0b1(din_26_ab1), .a0b2(din_26_ab2), .a0b3(din_26_ab3),
           .a0b0_1sc(din_26_ab0_1sc), .a0b1_1sc(din_26_ab1_1sc), .a0b2_1sc(din_26_ab2_1sc), .a0b3_1sc(din_26_ab3_1sc),
           .msk_a0b0(din_26_msk_ab0), .msk_a0b1(din_26_msk_ab1), .msk_a0b2(din_26_msk_ab2), .msk_a0b3(din_26_msk_ab3),
           .msk_a0b0_1sc(din_26_msk_ab0_1sc), .msk_a0b1_1sc(din_26_msk_ab1_1sc), .msk_a0b2_1sc(din_26_msk_ab2_1sc), .msk_a0b3_1sc(din_26_msk_ab3_1sc),

           .a1b0(din_28_ab0), .a1b1(din_28_ab1), .a1b2(din_28_ab2),
           .a1b0_1sc(din_28_ab0_1sc), .a1b1_1sc(din_28_ab1_1sc), .a1b2_1sc(din_28_ab2_1sc),
           .msk_a1b0(din_28_msk_ab0), .msk_a1b1(din_28_msk_ab1), .msk_a1b2(din_28_msk_ab2),
           .msk_a1b0_1sc(din_28_msk_ab0_1sc), .msk_a1b1_1sc(din_28_msk_ab1_1sc), .msk_a1b2_1sc(din_28_msk_ab2_1sc),

           .a2b0(din_30_ab0), .a2b1(din_30_ab1),
           .a2b0_1sc(din_30_ab0_1sc), .a2b1_1sc(din_30_ab1_1sc),
           .msk_a2b0(din_30_msk_ab0), .msk_a2b1(din_30_msk_ab1),
           .msk_a2b0_1sc(din_30_msk_ab0_1sc), .msk_a2b1_1sc(din_30_msk_ab1_1sc),
           
           .a3b0(din_32_ab0),
           .a3b0_1sc(din_32_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_27_calc (
           .clk(clk), .sign(din_signs_reg[27]), 
           .p(addr_3_27),
           .a0b0(din_27_ab0), .a0b1(din_27_ab1), .a0b2(din_27_ab2), .a0b3(din_27_ab3),
           .a0b0_1sc(din_27_ab0_1sc), .a0b1_1sc(din_27_ab1_1sc), .a0b2_1sc(din_27_ab2_1sc), .a0b3_1sc(din_27_ab3_1sc),
           .msk_a0b0(din_27_msk_ab0), .msk_a0b1(din_27_msk_ab1), .msk_a0b2(din_27_msk_ab2), .msk_a0b3(din_27_msk_ab3),
           .msk_a0b0_1sc(din_27_msk_ab0_1sc), .msk_a0b1_1sc(din_27_msk_ab1_1sc), .msk_a0b2_1sc(din_27_msk_ab2_1sc), .msk_a0b3_1sc(din_27_msk_ab3_1sc),

           .a1b0(din_29_ab0), .a1b1(din_29_ab1), .a1b2(din_29_ab2),
           .a1b0_1sc(din_29_ab0_1sc), .a1b1_1sc(din_29_ab1_1sc), .a1b2_1sc(din_29_ab2_1sc),
           .msk_a1b0(din_29_msk_ab0), .msk_a1b1(din_29_msk_ab1), .msk_a1b2(din_29_msk_ab2),
           .msk_a1b0_1sc(din_29_msk_ab0_1sc), .msk_a1b1_1sc(din_29_msk_ab1_1sc), .msk_a1b2_1sc(din_29_msk_ab2_1sc),

           .a2b0(din_31_ab0), .a2b1(din_31_ab1),
           .a2b0_1sc(din_31_ab0_1sc), .a2b1_1sc(din_31_ab1_1sc),
           .msk_a2b0(din_31_msk_ab0), .msk_a2b1(din_31_msk_ab1),
           .msk_a2b0_1sc(din_31_msk_ab0_1sc), .msk_a2b1_1sc(din_31_msk_ab1_1sc),
           
           .a3b0(din_33_ab0),
           .a3b0_1sc(din_33_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_28_calc (
           .clk(clk), .sign(din_signs_reg[28]), 
           .p(addr_3_28),
           .a0b0(din_28_ab0), .a0b1(din_28_ab1), .a0b2(din_28_ab2), .a0b3(din_28_ab3),
           .a0b0_1sc(din_28_ab0_1sc), .a0b1_1sc(din_28_ab1_1sc), .a0b2_1sc(din_28_ab2_1sc), .a0b3_1sc(din_28_ab3_1sc),
           .msk_a0b0(din_28_msk_ab0), .msk_a0b1(din_28_msk_ab1), .msk_a0b2(din_28_msk_ab2), .msk_a0b3(din_28_msk_ab3),
           .msk_a0b0_1sc(din_28_msk_ab0_1sc), .msk_a0b1_1sc(din_28_msk_ab1_1sc), .msk_a0b2_1sc(din_28_msk_ab2_1sc), .msk_a0b3_1sc(din_28_msk_ab3_1sc),

           .a1b0(din_30_ab0), .a1b1(din_30_ab1), .a1b2(din_30_ab2),
           .a1b0_1sc(din_30_ab0_1sc), .a1b1_1sc(din_30_ab1_1sc), .a1b2_1sc(din_30_ab2_1sc),
           .msk_a1b0(din_30_msk_ab0), .msk_a1b1(din_30_msk_ab1), .msk_a1b2(din_30_msk_ab2),
           .msk_a1b0_1sc(din_30_msk_ab0_1sc), .msk_a1b1_1sc(din_30_msk_ab1_1sc), .msk_a1b2_1sc(din_30_msk_ab2_1sc),

           .a2b0(din_32_ab0), .a2b1(din_32_ab1),
           .a2b0_1sc(din_32_ab0_1sc), .a2b1_1sc(din_32_ab1_1sc),
           .msk_a2b0(din_32_msk_ab0), .msk_a2b1(din_32_msk_ab1),
           .msk_a2b0_1sc(din_32_msk_ab0_1sc), .msk_a2b1_1sc(din_32_msk_ab1_1sc),
           
           .a3b0(din_34_ab0),
           .a3b0_1sc(din_34_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_29_calc (
           .clk(clk), .sign(din_signs_reg[29]), 
           .p(addr_3_29),
           .a0b0(din_29_ab0), .a0b1(din_29_ab1), .a0b2(din_29_ab2), .a0b3(din_29_ab3),
           .a0b0_1sc(din_29_ab0_1sc), .a0b1_1sc(din_29_ab1_1sc), .a0b2_1sc(din_29_ab2_1sc), .a0b3_1sc(din_29_ab3_1sc),
           .msk_a0b0(din_29_msk_ab0), .msk_a0b1(din_29_msk_ab1), .msk_a0b2(din_29_msk_ab2), .msk_a0b3(din_29_msk_ab3),
           .msk_a0b0_1sc(din_29_msk_ab0_1sc), .msk_a0b1_1sc(din_29_msk_ab1_1sc), .msk_a0b2_1sc(din_29_msk_ab2_1sc), .msk_a0b3_1sc(din_29_msk_ab3_1sc),

           .a1b0(din_31_ab0), .a1b1(din_31_ab1), .a1b2(din_31_ab2),
           .a1b0_1sc(din_31_ab0_1sc), .a1b1_1sc(din_31_ab1_1sc), .a1b2_1sc(din_31_ab2_1sc),
           .msk_a1b0(din_31_msk_ab0), .msk_a1b1(din_31_msk_ab1), .msk_a1b2(din_31_msk_ab2),
           .msk_a1b0_1sc(din_31_msk_ab0_1sc), .msk_a1b1_1sc(din_31_msk_ab1_1sc), .msk_a1b2_1sc(din_31_msk_ab2_1sc),

           .a2b0(din_33_ab0), .a2b1(din_33_ab1),
           .a2b0_1sc(din_33_ab0_1sc), .a2b1_1sc(din_33_ab1_1sc),
           .msk_a2b0(din_33_msk_ab0), .msk_a2b1(din_33_msk_ab1),
           .msk_a2b0_1sc(din_33_msk_ab0_1sc), .msk_a2b1_1sc(din_33_msk_ab1_1sc),
           
           .a3b0(din_35_ab0),
           .a3b0_1sc(din_35_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_30_calc (
           .clk(clk), .sign(din_signs_reg[30]), 
           .p(addr_3_30),
           .a0b0(din_30_ab0), .a0b1(din_30_ab1), .a0b2(din_30_ab2), .a0b3(din_30_ab3),
           .a0b0_1sc(din_30_ab0_1sc), .a0b1_1sc(din_30_ab1_1sc), .a0b2_1sc(din_30_ab2_1sc), .a0b3_1sc(din_30_ab3_1sc),
           .msk_a0b0(din_30_msk_ab0), .msk_a0b1(din_30_msk_ab1), .msk_a0b2(din_30_msk_ab2), .msk_a0b3(din_30_msk_ab3),
           .msk_a0b0_1sc(din_30_msk_ab0_1sc), .msk_a0b1_1sc(din_30_msk_ab1_1sc), .msk_a0b2_1sc(din_30_msk_ab2_1sc), .msk_a0b3_1sc(din_30_msk_ab3_1sc),

           .a1b0(din_32_ab0), .a1b1(din_32_ab1), .a1b2(din_32_ab2),
           .a1b0_1sc(din_32_ab0_1sc), .a1b1_1sc(din_32_ab1_1sc), .a1b2_1sc(din_32_ab2_1sc),
           .msk_a1b0(din_32_msk_ab0), .msk_a1b1(din_32_msk_ab1), .msk_a1b2(din_32_msk_ab2),
           .msk_a1b0_1sc(din_32_msk_ab0_1sc), .msk_a1b1_1sc(din_32_msk_ab1_1sc), .msk_a1b2_1sc(din_32_msk_ab2_1sc),

           .a2b0(din_34_ab0), .a2b1(din_34_ab1),
           .a2b0_1sc(din_34_ab0_1sc), .a2b1_1sc(din_34_ab1_1sc),
           .msk_a2b0(din_34_msk_ab0), .msk_a2b1(din_34_msk_ab1),
           .msk_a2b0_1sc(din_34_msk_ab0_1sc), .msk_a2b1_1sc(din_34_msk_ab1_1sc),
           
           .a3b0(din_36_ab0),
           .a3b0_1sc(din_36_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12)
) addr_3_31_calc (
           .clk(clk), .sign(din_signs_reg[31]), 
           .p(addr_3_31),
           .a0b0(din_31_ab0), .a0b1(din_31_ab1), .a0b2(din_31_ab2), .a0b3(din_31_ab3),
           .a0b0_1sc(din_31_ab0_1sc), .a0b1_1sc(din_31_ab1_1sc), .a0b2_1sc(din_31_ab2_1sc), .a0b3_1sc(din_31_ab3_1sc),
           .msk_a0b0(din_31_msk_ab0), .msk_a0b1(din_31_msk_ab1), .msk_a0b2(din_31_msk_ab2), .msk_a0b3(din_31_msk_ab3),
           .msk_a0b0_1sc(din_31_msk_ab0_1sc), .msk_a0b1_1sc(din_31_msk_ab1_1sc), .msk_a0b2_1sc(din_31_msk_ab2_1sc), .msk_a0b3_1sc(din_31_msk_ab3_1sc),

           .a1b0(din_33_ab0), .a1b1(din_33_ab1), .a1b2(din_33_ab2),
           .a1b0_1sc(din_33_ab0_1sc), .a1b1_1sc(din_33_ab1_1sc), .a1b2_1sc(din_33_ab2_1sc),
           .msk_a1b0(din_33_msk_ab0), .msk_a1b1(din_33_msk_ab1), .msk_a1b2(din_33_msk_ab2),
           .msk_a1b0_1sc(din_33_msk_ab0_1sc), .msk_a1b1_1sc(din_33_msk_ab1_1sc), .msk_a1b2_1sc(din_33_msk_ab2_1sc),

           .a2b0(din_35_ab0), .a2b1(din_35_ab1),
           .a2b0_1sc(din_35_ab0_1sc), .a2b1_1sc(din_35_ab1_1sc),
           .msk_a2b0(din_35_msk_ab0), .msk_a2b1(din_35_msk_ab1),
           .msk_a2b0_1sc(din_35_msk_ab0_1sc), .msk_a2b1_1sc(din_35_msk_ab1_1sc),
           
           .a3b0(din_37_ab0),
           .a3b0_1sc(din_37_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_0_calc (
           .clk(clk), .sign(din_signs_reg[0]), 
           .p(addr_4_0),
           .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
           .a0b0_1sc(din_0_ab0_1sc), .a0b1_1sc(din_0_ab1_1sc), .a0b2_1sc(din_0_ab2_1sc), .a0b3_1sc(din_0_ab3_1sc),
           .msk_a0b0(din_0_msk_ab0), .msk_a0b1(din_0_msk_ab1), .msk_a0b2(din_0_msk_ab2), .msk_a0b3(din_0_msk_ab3),
           .msk_a0b0_1sc(din_0_msk_ab0_1sc), .msk_a0b1_1sc(din_0_msk_ab1_1sc), .msk_a0b2_1sc(din_0_msk_ab2_1sc), .msk_a0b3_1sc(din_0_msk_ab3_1sc),

           .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2),
           .a1b0_1sc(din_2_ab0_1sc), .a1b1_1sc(din_2_ab1_1sc), .a1b2_1sc(din_2_ab2_1sc),
           .msk_a1b0(din_2_msk_ab0), .msk_a1b1(din_2_msk_ab1), .msk_a1b2(din_2_msk_ab2),
           .msk_a1b0_1sc(din_2_msk_ab0_1sc), .msk_a1b1_1sc(din_2_msk_ab1_1sc), .msk_a1b2_1sc(din_2_msk_ab2_1sc),

           .a2b0(din_4_ab0), .a2b1(din_4_ab1),
           .a2b0_1sc(din_4_ab0_1sc), .a2b1_1sc(din_4_ab1_1sc),
           .msk_a2b0(din_4_msk_ab0), .msk_a2b1(din_4_msk_ab1),
           .msk_a2b0_1sc(din_4_msk_ab0_1sc), .msk_a2b1_1sc(din_4_msk_ab1_1sc),
           
           .a3b0(din_6_ab0),
           .a3b0_1sc(din_6_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_1_calc (
           .clk(clk), .sign(din_signs_reg[1]), 
           .p(addr_4_1),
           .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
           .a0b0_1sc(din_1_ab0_1sc), .a0b1_1sc(din_1_ab1_1sc), .a0b2_1sc(din_1_ab2_1sc), .a0b3_1sc(din_1_ab3_1sc),
           .msk_a0b0(din_1_msk_ab0), .msk_a0b1(din_1_msk_ab1), .msk_a0b2(din_1_msk_ab2), .msk_a0b3(din_1_msk_ab3),
           .msk_a0b0_1sc(din_1_msk_ab0_1sc), .msk_a0b1_1sc(din_1_msk_ab1_1sc), .msk_a0b2_1sc(din_1_msk_ab2_1sc), .msk_a0b3_1sc(din_1_msk_ab3_1sc),

           .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2),
           .a1b0_1sc(din_3_ab0_1sc), .a1b1_1sc(din_3_ab1_1sc), .a1b2_1sc(din_3_ab2_1sc),
           .msk_a1b0(din_3_msk_ab0), .msk_a1b1(din_3_msk_ab1), .msk_a1b2(din_3_msk_ab2),
           .msk_a1b0_1sc(din_3_msk_ab0_1sc), .msk_a1b1_1sc(din_3_msk_ab1_1sc), .msk_a1b2_1sc(din_3_msk_ab2_1sc),

           .a2b0(din_5_ab0), .a2b1(din_5_ab1),
           .a2b0_1sc(din_5_ab0_1sc), .a2b1_1sc(din_5_ab1_1sc),
           .msk_a2b0(din_5_msk_ab0), .msk_a2b1(din_5_msk_ab1),
           .msk_a2b0_1sc(din_5_msk_ab0_1sc), .msk_a2b1_1sc(din_5_msk_ab1_1sc),
           
           .a3b0(din_7_ab0),
           .a3b0_1sc(din_7_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_2_calc (
           .clk(clk), .sign(din_signs_reg[2]), 
           .p(addr_4_2),
           .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
           .a0b0_1sc(din_2_ab0_1sc), .a0b1_1sc(din_2_ab1_1sc), .a0b2_1sc(din_2_ab2_1sc), .a0b3_1sc(din_2_ab3_1sc),
           .msk_a0b0(din_2_msk_ab0), .msk_a0b1(din_2_msk_ab1), .msk_a0b2(din_2_msk_ab2), .msk_a0b3(din_2_msk_ab3),
           .msk_a0b0_1sc(din_2_msk_ab0_1sc), .msk_a0b1_1sc(din_2_msk_ab1_1sc), .msk_a0b2_1sc(din_2_msk_ab2_1sc), .msk_a0b3_1sc(din_2_msk_ab3_1sc),

           .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2),
           .a1b0_1sc(din_4_ab0_1sc), .a1b1_1sc(din_4_ab1_1sc), .a1b2_1sc(din_4_ab2_1sc),
           .msk_a1b0(din_4_msk_ab0), .msk_a1b1(din_4_msk_ab1), .msk_a1b2(din_4_msk_ab2),
           .msk_a1b0_1sc(din_4_msk_ab0_1sc), .msk_a1b1_1sc(din_4_msk_ab1_1sc), .msk_a1b2_1sc(din_4_msk_ab2_1sc),

           .a2b0(din_6_ab0), .a2b1(din_6_ab1),
           .a2b0_1sc(din_6_ab0_1sc), .a2b1_1sc(din_6_ab1_1sc),
           .msk_a2b0(din_6_msk_ab0), .msk_a2b1(din_6_msk_ab1),
           .msk_a2b0_1sc(din_6_msk_ab0_1sc), .msk_a2b1_1sc(din_6_msk_ab1_1sc),
           
           .a3b0(din_8_ab0),
           .a3b0_1sc(din_8_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_3_calc (
           .clk(clk), .sign(din_signs_reg[3]), 
           .p(addr_4_3),
           .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
           .a0b0_1sc(din_3_ab0_1sc), .a0b1_1sc(din_3_ab1_1sc), .a0b2_1sc(din_3_ab2_1sc), .a0b3_1sc(din_3_ab3_1sc),
           .msk_a0b0(din_3_msk_ab0), .msk_a0b1(din_3_msk_ab1), .msk_a0b2(din_3_msk_ab2), .msk_a0b3(din_3_msk_ab3),
           .msk_a0b0_1sc(din_3_msk_ab0_1sc), .msk_a0b1_1sc(din_3_msk_ab1_1sc), .msk_a0b2_1sc(din_3_msk_ab2_1sc), .msk_a0b3_1sc(din_3_msk_ab3_1sc),

           .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2),
           .a1b0_1sc(din_5_ab0_1sc), .a1b1_1sc(din_5_ab1_1sc), .a1b2_1sc(din_5_ab2_1sc),
           .msk_a1b0(din_5_msk_ab0), .msk_a1b1(din_5_msk_ab1), .msk_a1b2(din_5_msk_ab2),
           .msk_a1b0_1sc(din_5_msk_ab0_1sc), .msk_a1b1_1sc(din_5_msk_ab1_1sc), .msk_a1b2_1sc(din_5_msk_ab2_1sc),

           .a2b0(din_7_ab0), .a2b1(din_7_ab1),
           .a2b0_1sc(din_7_ab0_1sc), .a2b1_1sc(din_7_ab1_1sc),
           .msk_a2b0(din_7_msk_ab0), .msk_a2b1(din_7_msk_ab1),
           .msk_a2b0_1sc(din_7_msk_ab0_1sc), .msk_a2b1_1sc(din_7_msk_ab1_1sc),
           
           .a3b0(din_9_ab0),
           .a3b0_1sc(din_9_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_4_calc (
           .clk(clk), .sign(din_signs_reg[4]), 
           .p(addr_4_4),
           .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
           .a0b0_1sc(din_4_ab0_1sc), .a0b1_1sc(din_4_ab1_1sc), .a0b2_1sc(din_4_ab2_1sc), .a0b3_1sc(din_4_ab3_1sc),
           .msk_a0b0(din_4_msk_ab0), .msk_a0b1(din_4_msk_ab1), .msk_a0b2(din_4_msk_ab2), .msk_a0b3(din_4_msk_ab3),
           .msk_a0b0_1sc(din_4_msk_ab0_1sc), .msk_a0b1_1sc(din_4_msk_ab1_1sc), .msk_a0b2_1sc(din_4_msk_ab2_1sc), .msk_a0b3_1sc(din_4_msk_ab3_1sc),

           .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2),
           .a1b0_1sc(din_6_ab0_1sc), .a1b1_1sc(din_6_ab1_1sc), .a1b2_1sc(din_6_ab2_1sc),
           .msk_a1b0(din_6_msk_ab0), .msk_a1b1(din_6_msk_ab1), .msk_a1b2(din_6_msk_ab2),
           .msk_a1b0_1sc(din_6_msk_ab0_1sc), .msk_a1b1_1sc(din_6_msk_ab1_1sc), .msk_a1b2_1sc(din_6_msk_ab2_1sc),

           .a2b0(din_8_ab0), .a2b1(din_8_ab1),
           .a2b0_1sc(din_8_ab0_1sc), .a2b1_1sc(din_8_ab1_1sc),
           .msk_a2b0(din_8_msk_ab0), .msk_a2b1(din_8_msk_ab1),
           .msk_a2b0_1sc(din_8_msk_ab0_1sc), .msk_a2b1_1sc(din_8_msk_ab1_1sc),
           
           .a3b0(din_10_ab0),
           .a3b0_1sc(din_10_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_5_calc (
           .clk(clk), .sign(din_signs_reg[5]), 
           .p(addr_4_5),
           .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
           .a0b0_1sc(din_5_ab0_1sc), .a0b1_1sc(din_5_ab1_1sc), .a0b2_1sc(din_5_ab2_1sc), .a0b3_1sc(din_5_ab3_1sc),
           .msk_a0b0(din_5_msk_ab0), .msk_a0b1(din_5_msk_ab1), .msk_a0b2(din_5_msk_ab2), .msk_a0b3(din_5_msk_ab3),
           .msk_a0b0_1sc(din_5_msk_ab0_1sc), .msk_a0b1_1sc(din_5_msk_ab1_1sc), .msk_a0b2_1sc(din_5_msk_ab2_1sc), .msk_a0b3_1sc(din_5_msk_ab3_1sc),

           .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2),
           .a1b0_1sc(din_7_ab0_1sc), .a1b1_1sc(din_7_ab1_1sc), .a1b2_1sc(din_7_ab2_1sc),
           .msk_a1b0(din_7_msk_ab0), .msk_a1b1(din_7_msk_ab1), .msk_a1b2(din_7_msk_ab2),
           .msk_a1b0_1sc(din_7_msk_ab0_1sc), .msk_a1b1_1sc(din_7_msk_ab1_1sc), .msk_a1b2_1sc(din_7_msk_ab2_1sc),

           .a2b0(din_9_ab0), .a2b1(din_9_ab1),
           .a2b0_1sc(din_9_ab0_1sc), .a2b1_1sc(din_9_ab1_1sc),
           .msk_a2b0(din_9_msk_ab0), .msk_a2b1(din_9_msk_ab1),
           .msk_a2b0_1sc(din_9_msk_ab0_1sc), .msk_a2b1_1sc(din_9_msk_ab1_1sc),
           
           .a3b0(din_11_ab0),
           .a3b0_1sc(din_11_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_6_calc (
           .clk(clk), .sign(din_signs_reg[6]), 
           .p(addr_4_6),
           .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
           .a0b0_1sc(din_6_ab0_1sc), .a0b1_1sc(din_6_ab1_1sc), .a0b2_1sc(din_6_ab2_1sc), .a0b3_1sc(din_6_ab3_1sc),
           .msk_a0b0(din_6_msk_ab0), .msk_a0b1(din_6_msk_ab1), .msk_a0b2(din_6_msk_ab2), .msk_a0b3(din_6_msk_ab3),
           .msk_a0b0_1sc(din_6_msk_ab0_1sc), .msk_a0b1_1sc(din_6_msk_ab1_1sc), .msk_a0b2_1sc(din_6_msk_ab2_1sc), .msk_a0b3_1sc(din_6_msk_ab3_1sc),

           .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2),
           .a1b0_1sc(din_8_ab0_1sc), .a1b1_1sc(din_8_ab1_1sc), .a1b2_1sc(din_8_ab2_1sc),
           .msk_a1b0(din_8_msk_ab0), .msk_a1b1(din_8_msk_ab1), .msk_a1b2(din_8_msk_ab2),
           .msk_a1b0_1sc(din_8_msk_ab0_1sc), .msk_a1b1_1sc(din_8_msk_ab1_1sc), .msk_a1b2_1sc(din_8_msk_ab2_1sc),

           .a2b0(din_10_ab0), .a2b1(din_10_ab1),
           .a2b0_1sc(din_10_ab0_1sc), .a2b1_1sc(din_10_ab1_1sc),
           .msk_a2b0(din_10_msk_ab0), .msk_a2b1(din_10_msk_ab1),
           .msk_a2b0_1sc(din_10_msk_ab0_1sc), .msk_a2b1_1sc(din_10_msk_ab1_1sc),
           
           .a3b0(din_12_ab0),
           .a3b0_1sc(din_12_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_7_calc (
           .clk(clk), .sign(din_signs_reg[7]), 
           .p(addr_4_7),
           .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
           .a0b0_1sc(din_7_ab0_1sc), .a0b1_1sc(din_7_ab1_1sc), .a0b2_1sc(din_7_ab2_1sc), .a0b3_1sc(din_7_ab3_1sc),
           .msk_a0b0(din_7_msk_ab0), .msk_a0b1(din_7_msk_ab1), .msk_a0b2(din_7_msk_ab2), .msk_a0b3(din_7_msk_ab3),
           .msk_a0b0_1sc(din_7_msk_ab0_1sc), .msk_a0b1_1sc(din_7_msk_ab1_1sc), .msk_a0b2_1sc(din_7_msk_ab2_1sc), .msk_a0b3_1sc(din_7_msk_ab3_1sc),

           .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2),
           .a1b0_1sc(din_9_ab0_1sc), .a1b1_1sc(din_9_ab1_1sc), .a1b2_1sc(din_9_ab2_1sc),
           .msk_a1b0(din_9_msk_ab0), .msk_a1b1(din_9_msk_ab1), .msk_a1b2(din_9_msk_ab2),
           .msk_a1b0_1sc(din_9_msk_ab0_1sc), .msk_a1b1_1sc(din_9_msk_ab1_1sc), .msk_a1b2_1sc(din_9_msk_ab2_1sc),

           .a2b0(din_11_ab0), .a2b1(din_11_ab1),
           .a2b0_1sc(din_11_ab0_1sc), .a2b1_1sc(din_11_ab1_1sc),
           .msk_a2b0(din_11_msk_ab0), .msk_a2b1(din_11_msk_ab1),
           .msk_a2b0_1sc(din_11_msk_ab0_1sc), .msk_a2b1_1sc(din_11_msk_ab1_1sc),
           
           .a3b0(din_13_ab0),
           .a3b0_1sc(din_13_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_8_calc (
           .clk(clk), .sign(din_signs_reg[8]), 
           .p(addr_4_8),
           .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
           .a0b0_1sc(din_8_ab0_1sc), .a0b1_1sc(din_8_ab1_1sc), .a0b2_1sc(din_8_ab2_1sc), .a0b3_1sc(din_8_ab3_1sc),
           .msk_a0b0(din_8_msk_ab0), .msk_a0b1(din_8_msk_ab1), .msk_a0b2(din_8_msk_ab2), .msk_a0b3(din_8_msk_ab3),
           .msk_a0b0_1sc(din_8_msk_ab0_1sc), .msk_a0b1_1sc(din_8_msk_ab1_1sc), .msk_a0b2_1sc(din_8_msk_ab2_1sc), .msk_a0b3_1sc(din_8_msk_ab3_1sc),

           .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2),
           .a1b0_1sc(din_10_ab0_1sc), .a1b1_1sc(din_10_ab1_1sc), .a1b2_1sc(din_10_ab2_1sc),
           .msk_a1b0(din_10_msk_ab0), .msk_a1b1(din_10_msk_ab1), .msk_a1b2(din_10_msk_ab2),
           .msk_a1b0_1sc(din_10_msk_ab0_1sc), .msk_a1b1_1sc(din_10_msk_ab1_1sc), .msk_a1b2_1sc(din_10_msk_ab2_1sc),

           .a2b0(din_12_ab0), .a2b1(din_12_ab1),
           .a2b0_1sc(din_12_ab0_1sc), .a2b1_1sc(din_12_ab1_1sc),
           .msk_a2b0(din_12_msk_ab0), .msk_a2b1(din_12_msk_ab1),
           .msk_a2b0_1sc(din_12_msk_ab0_1sc), .msk_a2b1_1sc(din_12_msk_ab1_1sc),
           
           .a3b0(din_14_ab0),
           .a3b0_1sc(din_14_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_9_calc (
           .clk(clk), .sign(din_signs_reg[9]), 
           .p(addr_4_9),
           .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
           .a0b0_1sc(din_9_ab0_1sc), .a0b1_1sc(din_9_ab1_1sc), .a0b2_1sc(din_9_ab2_1sc), .a0b3_1sc(din_9_ab3_1sc),
           .msk_a0b0(din_9_msk_ab0), .msk_a0b1(din_9_msk_ab1), .msk_a0b2(din_9_msk_ab2), .msk_a0b3(din_9_msk_ab3),
           .msk_a0b0_1sc(din_9_msk_ab0_1sc), .msk_a0b1_1sc(din_9_msk_ab1_1sc), .msk_a0b2_1sc(din_9_msk_ab2_1sc), .msk_a0b3_1sc(din_9_msk_ab3_1sc),

           .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2),
           .a1b0_1sc(din_11_ab0_1sc), .a1b1_1sc(din_11_ab1_1sc), .a1b2_1sc(din_11_ab2_1sc),
           .msk_a1b0(din_11_msk_ab0), .msk_a1b1(din_11_msk_ab1), .msk_a1b2(din_11_msk_ab2),
           .msk_a1b0_1sc(din_11_msk_ab0_1sc), .msk_a1b1_1sc(din_11_msk_ab1_1sc), .msk_a1b2_1sc(din_11_msk_ab2_1sc),

           .a2b0(din_13_ab0), .a2b1(din_13_ab1),
           .a2b0_1sc(din_13_ab0_1sc), .a2b1_1sc(din_13_ab1_1sc),
           .msk_a2b0(din_13_msk_ab0), .msk_a2b1(din_13_msk_ab1),
           .msk_a2b0_1sc(din_13_msk_ab0_1sc), .msk_a2b1_1sc(din_13_msk_ab1_1sc),
           
           .a3b0(din_15_ab0),
           .a3b0_1sc(din_15_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_10_calc (
           .clk(clk), .sign(din_signs_reg[10]), 
           .p(addr_4_10),
           .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
           .a0b0_1sc(din_10_ab0_1sc), .a0b1_1sc(din_10_ab1_1sc), .a0b2_1sc(din_10_ab2_1sc), .a0b3_1sc(din_10_ab3_1sc),
           .msk_a0b0(din_10_msk_ab0), .msk_a0b1(din_10_msk_ab1), .msk_a0b2(din_10_msk_ab2), .msk_a0b3(din_10_msk_ab3),
           .msk_a0b0_1sc(din_10_msk_ab0_1sc), .msk_a0b1_1sc(din_10_msk_ab1_1sc), .msk_a0b2_1sc(din_10_msk_ab2_1sc), .msk_a0b3_1sc(din_10_msk_ab3_1sc),

           .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2),
           .a1b0_1sc(din_12_ab0_1sc), .a1b1_1sc(din_12_ab1_1sc), .a1b2_1sc(din_12_ab2_1sc),
           .msk_a1b0(din_12_msk_ab0), .msk_a1b1(din_12_msk_ab1), .msk_a1b2(din_12_msk_ab2),
           .msk_a1b0_1sc(din_12_msk_ab0_1sc), .msk_a1b1_1sc(din_12_msk_ab1_1sc), .msk_a1b2_1sc(din_12_msk_ab2_1sc),

           .a2b0(din_14_ab0), .a2b1(din_14_ab1),
           .a2b0_1sc(din_14_ab0_1sc), .a2b1_1sc(din_14_ab1_1sc),
           .msk_a2b0(din_14_msk_ab0), .msk_a2b1(din_14_msk_ab1),
           .msk_a2b0_1sc(din_14_msk_ab0_1sc), .msk_a2b1_1sc(din_14_msk_ab1_1sc),
           
           .a3b0(din_16_ab0),
           .a3b0_1sc(din_16_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_11_calc (
           .clk(clk), .sign(din_signs_reg[11]), 
           .p(addr_4_11),
           .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
           .a0b0_1sc(din_11_ab0_1sc), .a0b1_1sc(din_11_ab1_1sc), .a0b2_1sc(din_11_ab2_1sc), .a0b3_1sc(din_11_ab3_1sc),
           .msk_a0b0(din_11_msk_ab0), .msk_a0b1(din_11_msk_ab1), .msk_a0b2(din_11_msk_ab2), .msk_a0b3(din_11_msk_ab3),
           .msk_a0b0_1sc(din_11_msk_ab0_1sc), .msk_a0b1_1sc(din_11_msk_ab1_1sc), .msk_a0b2_1sc(din_11_msk_ab2_1sc), .msk_a0b3_1sc(din_11_msk_ab3_1sc),

           .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2),
           .a1b0_1sc(din_13_ab0_1sc), .a1b1_1sc(din_13_ab1_1sc), .a1b2_1sc(din_13_ab2_1sc),
           .msk_a1b0(din_13_msk_ab0), .msk_a1b1(din_13_msk_ab1), .msk_a1b2(din_13_msk_ab2),
           .msk_a1b0_1sc(din_13_msk_ab0_1sc), .msk_a1b1_1sc(din_13_msk_ab1_1sc), .msk_a1b2_1sc(din_13_msk_ab2_1sc),

           .a2b0(din_15_ab0), .a2b1(din_15_ab1),
           .a2b0_1sc(din_15_ab0_1sc), .a2b1_1sc(din_15_ab1_1sc),
           .msk_a2b0(din_15_msk_ab0), .msk_a2b1(din_15_msk_ab1),
           .msk_a2b0_1sc(din_15_msk_ab0_1sc), .msk_a2b1_1sc(din_15_msk_ab1_1sc),
           
           .a3b0(din_17_ab0),
           .a3b0_1sc(din_17_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_12_calc (
           .clk(clk), .sign(din_signs_reg[12]), 
           .p(addr_4_12),
           .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
           .a0b0_1sc(din_12_ab0_1sc), .a0b1_1sc(din_12_ab1_1sc), .a0b2_1sc(din_12_ab2_1sc), .a0b3_1sc(din_12_ab3_1sc),
           .msk_a0b0(din_12_msk_ab0), .msk_a0b1(din_12_msk_ab1), .msk_a0b2(din_12_msk_ab2), .msk_a0b3(din_12_msk_ab3),
           .msk_a0b0_1sc(din_12_msk_ab0_1sc), .msk_a0b1_1sc(din_12_msk_ab1_1sc), .msk_a0b2_1sc(din_12_msk_ab2_1sc), .msk_a0b3_1sc(din_12_msk_ab3_1sc),

           .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2),
           .a1b0_1sc(din_14_ab0_1sc), .a1b1_1sc(din_14_ab1_1sc), .a1b2_1sc(din_14_ab2_1sc),
           .msk_a1b0(din_14_msk_ab0), .msk_a1b1(din_14_msk_ab1), .msk_a1b2(din_14_msk_ab2),
           .msk_a1b0_1sc(din_14_msk_ab0_1sc), .msk_a1b1_1sc(din_14_msk_ab1_1sc), .msk_a1b2_1sc(din_14_msk_ab2_1sc),

           .a2b0(din_16_ab0), .a2b1(din_16_ab1),
           .a2b0_1sc(din_16_ab0_1sc), .a2b1_1sc(din_16_ab1_1sc),
           .msk_a2b0(din_16_msk_ab0), .msk_a2b1(din_16_msk_ab1),
           .msk_a2b0_1sc(din_16_msk_ab0_1sc), .msk_a2b1_1sc(din_16_msk_ab1_1sc),
           
           .a3b0(din_18_ab0),
           .a3b0_1sc(din_18_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_13_calc (
           .clk(clk), .sign(din_signs_reg[13]), 
           .p(addr_4_13),
           .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
           .a0b0_1sc(din_13_ab0_1sc), .a0b1_1sc(din_13_ab1_1sc), .a0b2_1sc(din_13_ab2_1sc), .a0b3_1sc(din_13_ab3_1sc),
           .msk_a0b0(din_13_msk_ab0), .msk_a0b1(din_13_msk_ab1), .msk_a0b2(din_13_msk_ab2), .msk_a0b3(din_13_msk_ab3),
           .msk_a0b0_1sc(din_13_msk_ab0_1sc), .msk_a0b1_1sc(din_13_msk_ab1_1sc), .msk_a0b2_1sc(din_13_msk_ab2_1sc), .msk_a0b3_1sc(din_13_msk_ab3_1sc),

           .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2),
           .a1b0_1sc(din_15_ab0_1sc), .a1b1_1sc(din_15_ab1_1sc), .a1b2_1sc(din_15_ab2_1sc),
           .msk_a1b0(din_15_msk_ab0), .msk_a1b1(din_15_msk_ab1), .msk_a1b2(din_15_msk_ab2),
           .msk_a1b0_1sc(din_15_msk_ab0_1sc), .msk_a1b1_1sc(din_15_msk_ab1_1sc), .msk_a1b2_1sc(din_15_msk_ab2_1sc),

           .a2b0(din_17_ab0), .a2b1(din_17_ab1),
           .a2b0_1sc(din_17_ab0_1sc), .a2b1_1sc(din_17_ab1_1sc),
           .msk_a2b0(din_17_msk_ab0), .msk_a2b1(din_17_msk_ab1),
           .msk_a2b0_1sc(din_17_msk_ab0_1sc), .msk_a2b1_1sc(din_17_msk_ab1_1sc),
           
           .a3b0(din_19_ab0),
           .a3b0_1sc(din_19_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_14_calc (
           .clk(clk), .sign(din_signs_reg[14]), 
           .p(addr_4_14),
           .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
           .a0b0_1sc(din_14_ab0_1sc), .a0b1_1sc(din_14_ab1_1sc), .a0b2_1sc(din_14_ab2_1sc), .a0b3_1sc(din_14_ab3_1sc),
           .msk_a0b0(din_14_msk_ab0), .msk_a0b1(din_14_msk_ab1), .msk_a0b2(din_14_msk_ab2), .msk_a0b3(din_14_msk_ab3),
           .msk_a0b0_1sc(din_14_msk_ab0_1sc), .msk_a0b1_1sc(din_14_msk_ab1_1sc), .msk_a0b2_1sc(din_14_msk_ab2_1sc), .msk_a0b3_1sc(din_14_msk_ab3_1sc),

           .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2),
           .a1b0_1sc(din_16_ab0_1sc), .a1b1_1sc(din_16_ab1_1sc), .a1b2_1sc(din_16_ab2_1sc),
           .msk_a1b0(din_16_msk_ab0), .msk_a1b1(din_16_msk_ab1), .msk_a1b2(din_16_msk_ab2),
           .msk_a1b0_1sc(din_16_msk_ab0_1sc), .msk_a1b1_1sc(din_16_msk_ab1_1sc), .msk_a1b2_1sc(din_16_msk_ab2_1sc),

           .a2b0(din_18_ab0), .a2b1(din_18_ab1),
           .a2b0_1sc(din_18_ab0_1sc), .a2b1_1sc(din_18_ab1_1sc),
           .msk_a2b0(din_18_msk_ab0), .msk_a2b1(din_18_msk_ab1),
           .msk_a2b0_1sc(din_18_msk_ab0_1sc), .msk_a2b1_1sc(din_18_msk_ab1_1sc),
           
           .a3b0(din_20_ab0),
           .a3b0_1sc(din_20_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_15_calc (
           .clk(clk), .sign(din_signs_reg[15]), 
           .p(addr_4_15),
           .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
           .a0b0_1sc(din_15_ab0_1sc), .a0b1_1sc(din_15_ab1_1sc), .a0b2_1sc(din_15_ab2_1sc), .a0b3_1sc(din_15_ab3_1sc),
           .msk_a0b0(din_15_msk_ab0), .msk_a0b1(din_15_msk_ab1), .msk_a0b2(din_15_msk_ab2), .msk_a0b3(din_15_msk_ab3),
           .msk_a0b0_1sc(din_15_msk_ab0_1sc), .msk_a0b1_1sc(din_15_msk_ab1_1sc), .msk_a0b2_1sc(din_15_msk_ab2_1sc), .msk_a0b3_1sc(din_15_msk_ab3_1sc),

           .a1b0(din_17_ab0), .a1b1(din_17_ab1), .a1b2(din_17_ab2),
           .a1b0_1sc(din_17_ab0_1sc), .a1b1_1sc(din_17_ab1_1sc), .a1b2_1sc(din_17_ab2_1sc),
           .msk_a1b0(din_17_msk_ab0), .msk_a1b1(din_17_msk_ab1), .msk_a1b2(din_17_msk_ab2),
           .msk_a1b0_1sc(din_17_msk_ab0_1sc), .msk_a1b1_1sc(din_17_msk_ab1_1sc), .msk_a1b2_1sc(din_17_msk_ab2_1sc),

           .a2b0(din_19_ab0), .a2b1(din_19_ab1),
           .a2b0_1sc(din_19_ab0_1sc), .a2b1_1sc(din_19_ab1_1sc),
           .msk_a2b0(din_19_msk_ab0), .msk_a2b1(din_19_msk_ab1),
           .msk_a2b0_1sc(din_19_msk_ab0_1sc), .msk_a2b1_1sc(din_19_msk_ab1_1sc),
           
           .a3b0(din_21_ab0),
           .a3b0_1sc(din_21_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_16_calc (
           .clk(clk), .sign(din_signs_reg[16]), 
           .p(addr_4_16),
           .a0b0(din_16_ab0), .a0b1(din_16_ab1), .a0b2(din_16_ab2), .a0b3(din_16_ab3),
           .a0b0_1sc(din_16_ab0_1sc), .a0b1_1sc(din_16_ab1_1sc), .a0b2_1sc(din_16_ab2_1sc), .a0b3_1sc(din_16_ab3_1sc),
           .msk_a0b0(din_16_msk_ab0), .msk_a0b1(din_16_msk_ab1), .msk_a0b2(din_16_msk_ab2), .msk_a0b3(din_16_msk_ab3),
           .msk_a0b0_1sc(din_16_msk_ab0_1sc), .msk_a0b1_1sc(din_16_msk_ab1_1sc), .msk_a0b2_1sc(din_16_msk_ab2_1sc), .msk_a0b3_1sc(din_16_msk_ab3_1sc),

           .a1b0(din_18_ab0), .a1b1(din_18_ab1), .a1b2(din_18_ab2),
           .a1b0_1sc(din_18_ab0_1sc), .a1b1_1sc(din_18_ab1_1sc), .a1b2_1sc(din_18_ab2_1sc),
           .msk_a1b0(din_18_msk_ab0), .msk_a1b1(din_18_msk_ab1), .msk_a1b2(din_18_msk_ab2),
           .msk_a1b0_1sc(din_18_msk_ab0_1sc), .msk_a1b1_1sc(din_18_msk_ab1_1sc), .msk_a1b2_1sc(din_18_msk_ab2_1sc),

           .a2b0(din_20_ab0), .a2b1(din_20_ab1),
           .a2b0_1sc(din_20_ab0_1sc), .a2b1_1sc(din_20_ab1_1sc),
           .msk_a2b0(din_20_msk_ab0), .msk_a2b1(din_20_msk_ab1),
           .msk_a2b0_1sc(din_20_msk_ab0_1sc), .msk_a2b1_1sc(din_20_msk_ab1_1sc),
           
           .a3b0(din_22_ab0),
           .a3b0_1sc(din_22_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_17_calc (
           .clk(clk), .sign(din_signs_reg[17]), 
           .p(addr_4_17),
           .a0b0(din_17_ab0), .a0b1(din_17_ab1), .a0b2(din_17_ab2), .a0b3(din_17_ab3),
           .a0b0_1sc(din_17_ab0_1sc), .a0b1_1sc(din_17_ab1_1sc), .a0b2_1sc(din_17_ab2_1sc), .a0b3_1sc(din_17_ab3_1sc),
           .msk_a0b0(din_17_msk_ab0), .msk_a0b1(din_17_msk_ab1), .msk_a0b2(din_17_msk_ab2), .msk_a0b3(din_17_msk_ab3),
           .msk_a0b0_1sc(din_17_msk_ab0_1sc), .msk_a0b1_1sc(din_17_msk_ab1_1sc), .msk_a0b2_1sc(din_17_msk_ab2_1sc), .msk_a0b3_1sc(din_17_msk_ab3_1sc),

           .a1b0(din_19_ab0), .a1b1(din_19_ab1), .a1b2(din_19_ab2),
           .a1b0_1sc(din_19_ab0_1sc), .a1b1_1sc(din_19_ab1_1sc), .a1b2_1sc(din_19_ab2_1sc),
           .msk_a1b0(din_19_msk_ab0), .msk_a1b1(din_19_msk_ab1), .msk_a1b2(din_19_msk_ab2),
           .msk_a1b0_1sc(din_19_msk_ab0_1sc), .msk_a1b1_1sc(din_19_msk_ab1_1sc), .msk_a1b2_1sc(din_19_msk_ab2_1sc),

           .a2b0(din_21_ab0), .a2b1(din_21_ab1),
           .a2b0_1sc(din_21_ab0_1sc), .a2b1_1sc(din_21_ab1_1sc),
           .msk_a2b0(din_21_msk_ab0), .msk_a2b1(din_21_msk_ab1),
           .msk_a2b0_1sc(din_21_msk_ab0_1sc), .msk_a2b1_1sc(din_21_msk_ab1_1sc),
           
           .a3b0(din_23_ab0),
           .a3b0_1sc(din_23_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_18_calc (
           .clk(clk), .sign(din_signs_reg[18]), 
           .p(addr_4_18),
           .a0b0(din_18_ab0), .a0b1(din_18_ab1), .a0b2(din_18_ab2), .a0b3(din_18_ab3),
           .a0b0_1sc(din_18_ab0_1sc), .a0b1_1sc(din_18_ab1_1sc), .a0b2_1sc(din_18_ab2_1sc), .a0b3_1sc(din_18_ab3_1sc),
           .msk_a0b0(din_18_msk_ab0), .msk_a0b1(din_18_msk_ab1), .msk_a0b2(din_18_msk_ab2), .msk_a0b3(din_18_msk_ab3),
           .msk_a0b0_1sc(din_18_msk_ab0_1sc), .msk_a0b1_1sc(din_18_msk_ab1_1sc), .msk_a0b2_1sc(din_18_msk_ab2_1sc), .msk_a0b3_1sc(din_18_msk_ab3_1sc),

           .a1b0(din_20_ab0), .a1b1(din_20_ab1), .a1b2(din_20_ab2),
           .a1b0_1sc(din_20_ab0_1sc), .a1b1_1sc(din_20_ab1_1sc), .a1b2_1sc(din_20_ab2_1sc),
           .msk_a1b0(din_20_msk_ab0), .msk_a1b1(din_20_msk_ab1), .msk_a1b2(din_20_msk_ab2),
           .msk_a1b0_1sc(din_20_msk_ab0_1sc), .msk_a1b1_1sc(din_20_msk_ab1_1sc), .msk_a1b2_1sc(din_20_msk_ab2_1sc),

           .a2b0(din_22_ab0), .a2b1(din_22_ab1),
           .a2b0_1sc(din_22_ab0_1sc), .a2b1_1sc(din_22_ab1_1sc),
           .msk_a2b0(din_22_msk_ab0), .msk_a2b1(din_22_msk_ab1),
           .msk_a2b0_1sc(din_22_msk_ab0_1sc), .msk_a2b1_1sc(din_22_msk_ab1_1sc),
           
           .a3b0(din_24_ab0),
           .a3b0_1sc(din_24_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_19_calc (
           .clk(clk), .sign(din_signs_reg[19]), 
           .p(addr_4_19),
           .a0b0(din_19_ab0), .a0b1(din_19_ab1), .a0b2(din_19_ab2), .a0b3(din_19_ab3),
           .a0b0_1sc(din_19_ab0_1sc), .a0b1_1sc(din_19_ab1_1sc), .a0b2_1sc(din_19_ab2_1sc), .a0b3_1sc(din_19_ab3_1sc),
           .msk_a0b0(din_19_msk_ab0), .msk_a0b1(din_19_msk_ab1), .msk_a0b2(din_19_msk_ab2), .msk_a0b3(din_19_msk_ab3),
           .msk_a0b0_1sc(din_19_msk_ab0_1sc), .msk_a0b1_1sc(din_19_msk_ab1_1sc), .msk_a0b2_1sc(din_19_msk_ab2_1sc), .msk_a0b3_1sc(din_19_msk_ab3_1sc),

           .a1b0(din_21_ab0), .a1b1(din_21_ab1), .a1b2(din_21_ab2),
           .a1b0_1sc(din_21_ab0_1sc), .a1b1_1sc(din_21_ab1_1sc), .a1b2_1sc(din_21_ab2_1sc),
           .msk_a1b0(din_21_msk_ab0), .msk_a1b1(din_21_msk_ab1), .msk_a1b2(din_21_msk_ab2),
           .msk_a1b0_1sc(din_21_msk_ab0_1sc), .msk_a1b1_1sc(din_21_msk_ab1_1sc), .msk_a1b2_1sc(din_21_msk_ab2_1sc),

           .a2b0(din_23_ab0), .a2b1(din_23_ab1),
           .a2b0_1sc(din_23_ab0_1sc), .a2b1_1sc(din_23_ab1_1sc),
           .msk_a2b0(din_23_msk_ab0), .msk_a2b1(din_23_msk_ab1),
           .msk_a2b0_1sc(din_23_msk_ab0_1sc), .msk_a2b1_1sc(din_23_msk_ab1_1sc),
           
           .a3b0(din_25_ab0),
           .a3b0_1sc(din_25_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_20_calc (
           .clk(clk), .sign(din_signs_reg[20]), 
           .p(addr_4_20),
           .a0b0(din_20_ab0), .a0b1(din_20_ab1), .a0b2(din_20_ab2), .a0b3(din_20_ab3),
           .a0b0_1sc(din_20_ab0_1sc), .a0b1_1sc(din_20_ab1_1sc), .a0b2_1sc(din_20_ab2_1sc), .a0b3_1sc(din_20_ab3_1sc),
           .msk_a0b0(din_20_msk_ab0), .msk_a0b1(din_20_msk_ab1), .msk_a0b2(din_20_msk_ab2), .msk_a0b3(din_20_msk_ab3),
           .msk_a0b0_1sc(din_20_msk_ab0_1sc), .msk_a0b1_1sc(din_20_msk_ab1_1sc), .msk_a0b2_1sc(din_20_msk_ab2_1sc), .msk_a0b3_1sc(din_20_msk_ab3_1sc),

           .a1b0(din_22_ab0), .a1b1(din_22_ab1), .a1b2(din_22_ab2),
           .a1b0_1sc(din_22_ab0_1sc), .a1b1_1sc(din_22_ab1_1sc), .a1b2_1sc(din_22_ab2_1sc),
           .msk_a1b0(din_22_msk_ab0), .msk_a1b1(din_22_msk_ab1), .msk_a1b2(din_22_msk_ab2),
           .msk_a1b0_1sc(din_22_msk_ab0_1sc), .msk_a1b1_1sc(din_22_msk_ab1_1sc), .msk_a1b2_1sc(din_22_msk_ab2_1sc),

           .a2b0(din_24_ab0), .a2b1(din_24_ab1),
           .a2b0_1sc(din_24_ab0_1sc), .a2b1_1sc(din_24_ab1_1sc),
           .msk_a2b0(din_24_msk_ab0), .msk_a2b1(din_24_msk_ab1),
           .msk_a2b0_1sc(din_24_msk_ab0_1sc), .msk_a2b1_1sc(din_24_msk_ab1_1sc),
           
           .a3b0(din_26_ab0),
           .a3b0_1sc(din_26_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_21_calc (
           .clk(clk), .sign(din_signs_reg[21]), 
           .p(addr_4_21),
           .a0b0(din_21_ab0), .a0b1(din_21_ab1), .a0b2(din_21_ab2), .a0b3(din_21_ab3),
           .a0b0_1sc(din_21_ab0_1sc), .a0b1_1sc(din_21_ab1_1sc), .a0b2_1sc(din_21_ab2_1sc), .a0b3_1sc(din_21_ab3_1sc),
           .msk_a0b0(din_21_msk_ab0), .msk_a0b1(din_21_msk_ab1), .msk_a0b2(din_21_msk_ab2), .msk_a0b3(din_21_msk_ab3),
           .msk_a0b0_1sc(din_21_msk_ab0_1sc), .msk_a0b1_1sc(din_21_msk_ab1_1sc), .msk_a0b2_1sc(din_21_msk_ab2_1sc), .msk_a0b3_1sc(din_21_msk_ab3_1sc),

           .a1b0(din_23_ab0), .a1b1(din_23_ab1), .a1b2(din_23_ab2),
           .a1b0_1sc(din_23_ab0_1sc), .a1b1_1sc(din_23_ab1_1sc), .a1b2_1sc(din_23_ab2_1sc),
           .msk_a1b0(din_23_msk_ab0), .msk_a1b1(din_23_msk_ab1), .msk_a1b2(din_23_msk_ab2),
           .msk_a1b0_1sc(din_23_msk_ab0_1sc), .msk_a1b1_1sc(din_23_msk_ab1_1sc), .msk_a1b2_1sc(din_23_msk_ab2_1sc),

           .a2b0(din_25_ab0), .a2b1(din_25_ab1),
           .a2b0_1sc(din_25_ab0_1sc), .a2b1_1sc(din_25_ab1_1sc),
           .msk_a2b0(din_25_msk_ab0), .msk_a2b1(din_25_msk_ab1),
           .msk_a2b0_1sc(din_25_msk_ab0_1sc), .msk_a2b1_1sc(din_25_msk_ab1_1sc),
           
           .a3b0(din_27_ab0),
           .a3b0_1sc(din_27_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_22_calc (
           .clk(clk), .sign(din_signs_reg[22]), 
           .p(addr_4_22),
           .a0b0(din_22_ab0), .a0b1(din_22_ab1), .a0b2(din_22_ab2), .a0b3(din_22_ab3),
           .a0b0_1sc(din_22_ab0_1sc), .a0b1_1sc(din_22_ab1_1sc), .a0b2_1sc(din_22_ab2_1sc), .a0b3_1sc(din_22_ab3_1sc),
           .msk_a0b0(din_22_msk_ab0), .msk_a0b1(din_22_msk_ab1), .msk_a0b2(din_22_msk_ab2), .msk_a0b3(din_22_msk_ab3),
           .msk_a0b0_1sc(din_22_msk_ab0_1sc), .msk_a0b1_1sc(din_22_msk_ab1_1sc), .msk_a0b2_1sc(din_22_msk_ab2_1sc), .msk_a0b3_1sc(din_22_msk_ab3_1sc),

           .a1b0(din_24_ab0), .a1b1(din_24_ab1), .a1b2(din_24_ab2),
           .a1b0_1sc(din_24_ab0_1sc), .a1b1_1sc(din_24_ab1_1sc), .a1b2_1sc(din_24_ab2_1sc),
           .msk_a1b0(din_24_msk_ab0), .msk_a1b1(din_24_msk_ab1), .msk_a1b2(din_24_msk_ab2),
           .msk_a1b0_1sc(din_24_msk_ab0_1sc), .msk_a1b1_1sc(din_24_msk_ab1_1sc), .msk_a1b2_1sc(din_24_msk_ab2_1sc),

           .a2b0(din_26_ab0), .a2b1(din_26_ab1),
           .a2b0_1sc(din_26_ab0_1sc), .a2b1_1sc(din_26_ab1_1sc),
           .msk_a2b0(din_26_msk_ab0), .msk_a2b1(din_26_msk_ab1),
           .msk_a2b0_1sc(din_26_msk_ab0_1sc), .msk_a2b1_1sc(din_26_msk_ab1_1sc),
           
           .a3b0(din_28_ab0),
           .a3b0_1sc(din_28_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_23_calc (
           .clk(clk), .sign(din_signs_reg[23]), 
           .p(addr_4_23),
           .a0b0(din_23_ab0), .a0b1(din_23_ab1), .a0b2(din_23_ab2), .a0b3(din_23_ab3),
           .a0b0_1sc(din_23_ab0_1sc), .a0b1_1sc(din_23_ab1_1sc), .a0b2_1sc(din_23_ab2_1sc), .a0b3_1sc(din_23_ab3_1sc),
           .msk_a0b0(din_23_msk_ab0), .msk_a0b1(din_23_msk_ab1), .msk_a0b2(din_23_msk_ab2), .msk_a0b3(din_23_msk_ab3),
           .msk_a0b0_1sc(din_23_msk_ab0_1sc), .msk_a0b1_1sc(din_23_msk_ab1_1sc), .msk_a0b2_1sc(din_23_msk_ab2_1sc), .msk_a0b3_1sc(din_23_msk_ab3_1sc),

           .a1b0(din_25_ab0), .a1b1(din_25_ab1), .a1b2(din_25_ab2),
           .a1b0_1sc(din_25_ab0_1sc), .a1b1_1sc(din_25_ab1_1sc), .a1b2_1sc(din_25_ab2_1sc),
           .msk_a1b0(din_25_msk_ab0), .msk_a1b1(din_25_msk_ab1), .msk_a1b2(din_25_msk_ab2),
           .msk_a1b0_1sc(din_25_msk_ab0_1sc), .msk_a1b1_1sc(din_25_msk_ab1_1sc), .msk_a1b2_1sc(din_25_msk_ab2_1sc),

           .a2b0(din_27_ab0), .a2b1(din_27_ab1),
           .a2b0_1sc(din_27_ab0_1sc), .a2b1_1sc(din_27_ab1_1sc),
           .msk_a2b0(din_27_msk_ab0), .msk_a2b1(din_27_msk_ab1),
           .msk_a2b0_1sc(din_27_msk_ab0_1sc), .msk_a2b1_1sc(din_27_msk_ab1_1sc),
           
           .a3b0(din_29_ab0),
           .a3b0_1sc(din_29_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_24_calc (
           .clk(clk), .sign(din_signs_reg[24]), 
           .p(addr_4_24),
           .a0b0(din_24_ab0), .a0b1(din_24_ab1), .a0b2(din_24_ab2), .a0b3(din_24_ab3),
           .a0b0_1sc(din_24_ab0_1sc), .a0b1_1sc(din_24_ab1_1sc), .a0b2_1sc(din_24_ab2_1sc), .a0b3_1sc(din_24_ab3_1sc),
           .msk_a0b0(din_24_msk_ab0), .msk_a0b1(din_24_msk_ab1), .msk_a0b2(din_24_msk_ab2), .msk_a0b3(din_24_msk_ab3),
           .msk_a0b0_1sc(din_24_msk_ab0_1sc), .msk_a0b1_1sc(din_24_msk_ab1_1sc), .msk_a0b2_1sc(din_24_msk_ab2_1sc), .msk_a0b3_1sc(din_24_msk_ab3_1sc),

           .a1b0(din_26_ab0), .a1b1(din_26_ab1), .a1b2(din_26_ab2),
           .a1b0_1sc(din_26_ab0_1sc), .a1b1_1sc(din_26_ab1_1sc), .a1b2_1sc(din_26_ab2_1sc),
           .msk_a1b0(din_26_msk_ab0), .msk_a1b1(din_26_msk_ab1), .msk_a1b2(din_26_msk_ab2),
           .msk_a1b0_1sc(din_26_msk_ab0_1sc), .msk_a1b1_1sc(din_26_msk_ab1_1sc), .msk_a1b2_1sc(din_26_msk_ab2_1sc),

           .a2b0(din_28_ab0), .a2b1(din_28_ab1),
           .a2b0_1sc(din_28_ab0_1sc), .a2b1_1sc(din_28_ab1_1sc),
           .msk_a2b0(din_28_msk_ab0), .msk_a2b1(din_28_msk_ab1),
           .msk_a2b0_1sc(din_28_msk_ab0_1sc), .msk_a2b1_1sc(din_28_msk_ab1_1sc),
           
           .a3b0(din_30_ab0),
           .a3b0_1sc(din_30_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_25_calc (
           .clk(clk), .sign(din_signs_reg[25]), 
           .p(addr_4_25),
           .a0b0(din_25_ab0), .a0b1(din_25_ab1), .a0b2(din_25_ab2), .a0b3(din_25_ab3),
           .a0b0_1sc(din_25_ab0_1sc), .a0b1_1sc(din_25_ab1_1sc), .a0b2_1sc(din_25_ab2_1sc), .a0b3_1sc(din_25_ab3_1sc),
           .msk_a0b0(din_25_msk_ab0), .msk_a0b1(din_25_msk_ab1), .msk_a0b2(din_25_msk_ab2), .msk_a0b3(din_25_msk_ab3),
           .msk_a0b0_1sc(din_25_msk_ab0_1sc), .msk_a0b1_1sc(din_25_msk_ab1_1sc), .msk_a0b2_1sc(din_25_msk_ab2_1sc), .msk_a0b3_1sc(din_25_msk_ab3_1sc),

           .a1b0(din_27_ab0), .a1b1(din_27_ab1), .a1b2(din_27_ab2),
           .a1b0_1sc(din_27_ab0_1sc), .a1b1_1sc(din_27_ab1_1sc), .a1b2_1sc(din_27_ab2_1sc),
           .msk_a1b0(din_27_msk_ab0), .msk_a1b1(din_27_msk_ab1), .msk_a1b2(din_27_msk_ab2),
           .msk_a1b0_1sc(din_27_msk_ab0_1sc), .msk_a1b1_1sc(din_27_msk_ab1_1sc), .msk_a1b2_1sc(din_27_msk_ab2_1sc),

           .a2b0(din_29_ab0), .a2b1(din_29_ab1),
           .a2b0_1sc(din_29_ab0_1sc), .a2b1_1sc(din_29_ab1_1sc),
           .msk_a2b0(din_29_msk_ab0), .msk_a2b1(din_29_msk_ab1),
           .msk_a2b0_1sc(din_29_msk_ab0_1sc), .msk_a2b1_1sc(din_29_msk_ab1_1sc),
           
           .a3b0(din_31_ab0),
           .a3b0_1sc(din_31_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_26_calc (
           .clk(clk), .sign(din_signs_reg[26]), 
           .p(addr_4_26),
           .a0b0(din_26_ab0), .a0b1(din_26_ab1), .a0b2(din_26_ab2), .a0b3(din_26_ab3),
           .a0b0_1sc(din_26_ab0_1sc), .a0b1_1sc(din_26_ab1_1sc), .a0b2_1sc(din_26_ab2_1sc), .a0b3_1sc(din_26_ab3_1sc),
           .msk_a0b0(din_26_msk_ab0), .msk_a0b1(din_26_msk_ab1), .msk_a0b2(din_26_msk_ab2), .msk_a0b3(din_26_msk_ab3),
           .msk_a0b0_1sc(din_26_msk_ab0_1sc), .msk_a0b1_1sc(din_26_msk_ab1_1sc), .msk_a0b2_1sc(din_26_msk_ab2_1sc), .msk_a0b3_1sc(din_26_msk_ab3_1sc),

           .a1b0(din_28_ab0), .a1b1(din_28_ab1), .a1b2(din_28_ab2),
           .a1b0_1sc(din_28_ab0_1sc), .a1b1_1sc(din_28_ab1_1sc), .a1b2_1sc(din_28_ab2_1sc),
           .msk_a1b0(din_28_msk_ab0), .msk_a1b1(din_28_msk_ab1), .msk_a1b2(din_28_msk_ab2),
           .msk_a1b0_1sc(din_28_msk_ab0_1sc), .msk_a1b1_1sc(din_28_msk_ab1_1sc), .msk_a1b2_1sc(din_28_msk_ab2_1sc),

           .a2b0(din_30_ab0), .a2b1(din_30_ab1),
           .a2b0_1sc(din_30_ab0_1sc), .a2b1_1sc(din_30_ab1_1sc),
           .msk_a2b0(din_30_msk_ab0), .msk_a2b1(din_30_msk_ab1),
           .msk_a2b0_1sc(din_30_msk_ab0_1sc), .msk_a2b1_1sc(din_30_msk_ab1_1sc),
           
           .a3b0(din_32_ab0),
           .a3b0_1sc(din_32_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_27_calc (
           .clk(clk), .sign(din_signs_reg[27]), 
           .p(addr_4_27),
           .a0b0(din_27_ab0), .a0b1(din_27_ab1), .a0b2(din_27_ab2), .a0b3(din_27_ab3),
           .a0b0_1sc(din_27_ab0_1sc), .a0b1_1sc(din_27_ab1_1sc), .a0b2_1sc(din_27_ab2_1sc), .a0b3_1sc(din_27_ab3_1sc),
           .msk_a0b0(din_27_msk_ab0), .msk_a0b1(din_27_msk_ab1), .msk_a0b2(din_27_msk_ab2), .msk_a0b3(din_27_msk_ab3),
           .msk_a0b0_1sc(din_27_msk_ab0_1sc), .msk_a0b1_1sc(din_27_msk_ab1_1sc), .msk_a0b2_1sc(din_27_msk_ab2_1sc), .msk_a0b3_1sc(din_27_msk_ab3_1sc),

           .a1b0(din_29_ab0), .a1b1(din_29_ab1), .a1b2(din_29_ab2),
           .a1b0_1sc(din_29_ab0_1sc), .a1b1_1sc(din_29_ab1_1sc), .a1b2_1sc(din_29_ab2_1sc),
           .msk_a1b0(din_29_msk_ab0), .msk_a1b1(din_29_msk_ab1), .msk_a1b2(din_29_msk_ab2),
           .msk_a1b0_1sc(din_29_msk_ab0_1sc), .msk_a1b1_1sc(din_29_msk_ab1_1sc), .msk_a1b2_1sc(din_29_msk_ab2_1sc),

           .a2b0(din_31_ab0), .a2b1(din_31_ab1),
           .a2b0_1sc(din_31_ab0_1sc), .a2b1_1sc(din_31_ab1_1sc),
           .msk_a2b0(din_31_msk_ab0), .msk_a2b1(din_31_msk_ab1),
           .msk_a2b0_1sc(din_31_msk_ab0_1sc), .msk_a2b1_1sc(din_31_msk_ab1_1sc),
           
           .a3b0(din_33_ab0),
           .a3b0_1sc(din_33_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_28_calc (
           .clk(clk), .sign(din_signs_reg[28]), 
           .p(addr_4_28),
           .a0b0(din_28_ab0), .a0b1(din_28_ab1), .a0b2(din_28_ab2), .a0b3(din_28_ab3),
           .a0b0_1sc(din_28_ab0_1sc), .a0b1_1sc(din_28_ab1_1sc), .a0b2_1sc(din_28_ab2_1sc), .a0b3_1sc(din_28_ab3_1sc),
           .msk_a0b0(din_28_msk_ab0), .msk_a0b1(din_28_msk_ab1), .msk_a0b2(din_28_msk_ab2), .msk_a0b3(din_28_msk_ab3),
           .msk_a0b0_1sc(din_28_msk_ab0_1sc), .msk_a0b1_1sc(din_28_msk_ab1_1sc), .msk_a0b2_1sc(din_28_msk_ab2_1sc), .msk_a0b3_1sc(din_28_msk_ab3_1sc),

           .a1b0(din_30_ab0), .a1b1(din_30_ab1), .a1b2(din_30_ab2),
           .a1b0_1sc(din_30_ab0_1sc), .a1b1_1sc(din_30_ab1_1sc), .a1b2_1sc(din_30_ab2_1sc),
           .msk_a1b0(din_30_msk_ab0), .msk_a1b1(din_30_msk_ab1), .msk_a1b2(din_30_msk_ab2),
           .msk_a1b0_1sc(din_30_msk_ab0_1sc), .msk_a1b1_1sc(din_30_msk_ab1_1sc), .msk_a1b2_1sc(din_30_msk_ab2_1sc),

           .a2b0(din_32_ab0), .a2b1(din_32_ab1),
           .a2b0_1sc(din_32_ab0_1sc), .a2b1_1sc(din_32_ab1_1sc),
           .msk_a2b0(din_32_msk_ab0), .msk_a2b1(din_32_msk_ab1),
           .msk_a2b0_1sc(din_32_msk_ab0_1sc), .msk_a2b1_1sc(din_32_msk_ab1_1sc),
           
           .a3b0(din_34_ab0),
           .a3b0_1sc(din_34_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_29_calc (
           .clk(clk), .sign(din_signs_reg[29]), 
           .p(addr_4_29),
           .a0b0(din_29_ab0), .a0b1(din_29_ab1), .a0b2(din_29_ab2), .a0b3(din_29_ab3),
           .a0b0_1sc(din_29_ab0_1sc), .a0b1_1sc(din_29_ab1_1sc), .a0b2_1sc(din_29_ab2_1sc), .a0b3_1sc(din_29_ab3_1sc),
           .msk_a0b0(din_29_msk_ab0), .msk_a0b1(din_29_msk_ab1), .msk_a0b2(din_29_msk_ab2), .msk_a0b3(din_29_msk_ab3),
           .msk_a0b0_1sc(din_29_msk_ab0_1sc), .msk_a0b1_1sc(din_29_msk_ab1_1sc), .msk_a0b2_1sc(din_29_msk_ab2_1sc), .msk_a0b3_1sc(din_29_msk_ab3_1sc),

           .a1b0(din_31_ab0), .a1b1(din_31_ab1), .a1b2(din_31_ab2),
           .a1b0_1sc(din_31_ab0_1sc), .a1b1_1sc(din_31_ab1_1sc), .a1b2_1sc(din_31_ab2_1sc),
           .msk_a1b0(din_31_msk_ab0), .msk_a1b1(din_31_msk_ab1), .msk_a1b2(din_31_msk_ab2),
           .msk_a1b0_1sc(din_31_msk_ab0_1sc), .msk_a1b1_1sc(din_31_msk_ab1_1sc), .msk_a1b2_1sc(din_31_msk_ab2_1sc),

           .a2b0(din_33_ab0), .a2b1(din_33_ab1),
           .a2b0_1sc(din_33_ab0_1sc), .a2b1_1sc(din_33_ab1_1sc),
           .msk_a2b0(din_33_msk_ab0), .msk_a2b1(din_33_msk_ab1),
           .msk_a2b0_1sc(din_33_msk_ab0_1sc), .msk_a2b1_1sc(din_33_msk_ab1_1sc),
           
           .a3b0(din_35_ab0),
           .a3b0_1sc(din_35_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_30_calc (
           .clk(clk), .sign(din_signs_reg[30]), 
           .p(addr_4_30),
           .a0b0(din_30_ab0), .a0b1(din_30_ab1), .a0b2(din_30_ab2), .a0b3(din_30_ab3),
           .a0b0_1sc(din_30_ab0_1sc), .a0b1_1sc(din_30_ab1_1sc), .a0b2_1sc(din_30_ab2_1sc), .a0b3_1sc(din_30_ab3_1sc),
           .msk_a0b0(din_30_msk_ab0), .msk_a0b1(din_30_msk_ab1), .msk_a0b2(din_30_msk_ab2), .msk_a0b3(din_30_msk_ab3),
           .msk_a0b0_1sc(din_30_msk_ab0_1sc), .msk_a0b1_1sc(din_30_msk_ab1_1sc), .msk_a0b2_1sc(din_30_msk_ab2_1sc), .msk_a0b3_1sc(din_30_msk_ab3_1sc),

           .a1b0(din_32_ab0), .a1b1(din_32_ab1), .a1b2(din_32_ab2),
           .a1b0_1sc(din_32_ab0_1sc), .a1b1_1sc(din_32_ab1_1sc), .a1b2_1sc(din_32_ab2_1sc),
           .msk_a1b0(din_32_msk_ab0), .msk_a1b1(din_32_msk_ab1), .msk_a1b2(din_32_msk_ab2),
           .msk_a1b0_1sc(din_32_msk_ab0_1sc), .msk_a1b1_1sc(din_32_msk_ab1_1sc), .msk_a1b2_1sc(din_32_msk_ab2_1sc),

           .a2b0(din_34_ab0), .a2b1(din_34_ab1),
           .a2b0_1sc(din_34_ab0_1sc), .a2b1_1sc(din_34_ab1_1sc),
           .msk_a2b0(din_34_msk_ab0), .msk_a2b1(din_34_msk_ab1),
           .msk_a2b0_1sc(din_34_msk_ab0_1sc), .msk_a2b1_1sc(din_34_msk_ab1_1sc),
           
           .a3b0(din_36_ab0),
           .a3b0_1sc(din_36_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11)
) addr_4_31_calc (
           .clk(clk), .sign(din_signs_reg[31]), 
           .p(addr_4_31),
           .a0b0(din_31_ab0), .a0b1(din_31_ab1), .a0b2(din_31_ab2), .a0b3(din_31_ab3),
           .a0b0_1sc(din_31_ab0_1sc), .a0b1_1sc(din_31_ab1_1sc), .a0b2_1sc(din_31_ab2_1sc), .a0b3_1sc(din_31_ab3_1sc),
           .msk_a0b0(din_31_msk_ab0), .msk_a0b1(din_31_msk_ab1), .msk_a0b2(din_31_msk_ab2), .msk_a0b3(din_31_msk_ab3),
           .msk_a0b0_1sc(din_31_msk_ab0_1sc), .msk_a0b1_1sc(din_31_msk_ab1_1sc), .msk_a0b2_1sc(din_31_msk_ab2_1sc), .msk_a0b3_1sc(din_31_msk_ab3_1sc),

           .a1b0(din_33_ab0), .a1b1(din_33_ab1), .a1b2(din_33_ab2),
           .a1b0_1sc(din_33_ab0_1sc), .a1b1_1sc(din_33_ab1_1sc), .a1b2_1sc(din_33_ab2_1sc),
           .msk_a1b0(din_33_msk_ab0), .msk_a1b1(din_33_msk_ab1), .msk_a1b2(din_33_msk_ab2),
           .msk_a1b0_1sc(din_33_msk_ab0_1sc), .msk_a1b1_1sc(din_33_msk_ab1_1sc), .msk_a1b2_1sc(din_33_msk_ab2_1sc),

           .a2b0(din_35_ab0), .a2b1(din_35_ab1),
           .a2b0_1sc(din_35_ab0_1sc), .a2b1_1sc(din_35_ab1_1sc),
           .msk_a2b0(din_35_msk_ab0), .msk_a2b1(din_35_msk_ab1),
           .msk_a2b0_1sc(din_35_msk_ab0_1sc), .msk_a2b1_1sc(din_35_msk_ab1_1sc),
           
           .a3b0(din_37_ab0),
           .a3b0_1sc(din_37_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_0_calc (
           .clk(clk), .sign(din_signs_reg[0]), 
           .p(addr_5_0),
           .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
           .a0b0_1sc(din_0_ab0_1sc), .a0b1_1sc(din_0_ab1_1sc), .a0b2_1sc(din_0_ab2_1sc), .a0b3_1sc(din_0_ab3_1sc),
           .msk_a0b0(din_0_msk_ab0), .msk_a0b1(din_0_msk_ab1), .msk_a0b2(din_0_msk_ab2), .msk_a0b3(din_0_msk_ab3),
           .msk_a0b0_1sc(din_0_msk_ab0_1sc), .msk_a0b1_1sc(din_0_msk_ab1_1sc), .msk_a0b2_1sc(din_0_msk_ab2_1sc), .msk_a0b3_1sc(din_0_msk_ab3_1sc),

           .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2),
           .a1b0_1sc(din_2_ab0_1sc), .a1b1_1sc(din_2_ab1_1sc), .a1b2_1sc(din_2_ab2_1sc),
           .msk_a1b0(din_2_msk_ab0), .msk_a1b1(din_2_msk_ab1), .msk_a1b2(din_2_msk_ab2),
           .msk_a1b0_1sc(din_2_msk_ab0_1sc), .msk_a1b1_1sc(din_2_msk_ab1_1sc), .msk_a1b2_1sc(din_2_msk_ab2_1sc),

           .a2b0(din_4_ab0), .a2b1(din_4_ab1),
           .a2b0_1sc(din_4_ab0_1sc), .a2b1_1sc(din_4_ab1_1sc),
           .msk_a2b0(din_4_msk_ab0), .msk_a2b1(din_4_msk_ab1),
           .msk_a2b0_1sc(din_4_msk_ab0_1sc), .msk_a2b1_1sc(din_4_msk_ab1_1sc),
           
           .a3b0(din_6_ab0),
           .a3b0_1sc(din_6_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_1_calc (
           .clk(clk), .sign(din_signs_reg[1]), 
           .p(addr_5_1),
           .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
           .a0b0_1sc(din_1_ab0_1sc), .a0b1_1sc(din_1_ab1_1sc), .a0b2_1sc(din_1_ab2_1sc), .a0b3_1sc(din_1_ab3_1sc),
           .msk_a0b0(din_1_msk_ab0), .msk_a0b1(din_1_msk_ab1), .msk_a0b2(din_1_msk_ab2), .msk_a0b3(din_1_msk_ab3),
           .msk_a0b0_1sc(din_1_msk_ab0_1sc), .msk_a0b1_1sc(din_1_msk_ab1_1sc), .msk_a0b2_1sc(din_1_msk_ab2_1sc), .msk_a0b3_1sc(din_1_msk_ab3_1sc),

           .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2),
           .a1b0_1sc(din_3_ab0_1sc), .a1b1_1sc(din_3_ab1_1sc), .a1b2_1sc(din_3_ab2_1sc),
           .msk_a1b0(din_3_msk_ab0), .msk_a1b1(din_3_msk_ab1), .msk_a1b2(din_3_msk_ab2),
           .msk_a1b0_1sc(din_3_msk_ab0_1sc), .msk_a1b1_1sc(din_3_msk_ab1_1sc), .msk_a1b2_1sc(din_3_msk_ab2_1sc),

           .a2b0(din_5_ab0), .a2b1(din_5_ab1),
           .a2b0_1sc(din_5_ab0_1sc), .a2b1_1sc(din_5_ab1_1sc),
           .msk_a2b0(din_5_msk_ab0), .msk_a2b1(din_5_msk_ab1),
           .msk_a2b0_1sc(din_5_msk_ab0_1sc), .msk_a2b1_1sc(din_5_msk_ab1_1sc),
           
           .a3b0(din_7_ab0),
           .a3b0_1sc(din_7_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_2_calc (
           .clk(clk), .sign(din_signs_reg[2]), 
           .p(addr_5_2),
           .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
           .a0b0_1sc(din_2_ab0_1sc), .a0b1_1sc(din_2_ab1_1sc), .a0b2_1sc(din_2_ab2_1sc), .a0b3_1sc(din_2_ab3_1sc),
           .msk_a0b0(din_2_msk_ab0), .msk_a0b1(din_2_msk_ab1), .msk_a0b2(din_2_msk_ab2), .msk_a0b3(din_2_msk_ab3),
           .msk_a0b0_1sc(din_2_msk_ab0_1sc), .msk_a0b1_1sc(din_2_msk_ab1_1sc), .msk_a0b2_1sc(din_2_msk_ab2_1sc), .msk_a0b3_1sc(din_2_msk_ab3_1sc),

           .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2),
           .a1b0_1sc(din_4_ab0_1sc), .a1b1_1sc(din_4_ab1_1sc), .a1b2_1sc(din_4_ab2_1sc),
           .msk_a1b0(din_4_msk_ab0), .msk_a1b1(din_4_msk_ab1), .msk_a1b2(din_4_msk_ab2),
           .msk_a1b0_1sc(din_4_msk_ab0_1sc), .msk_a1b1_1sc(din_4_msk_ab1_1sc), .msk_a1b2_1sc(din_4_msk_ab2_1sc),

           .a2b0(din_6_ab0), .a2b1(din_6_ab1),
           .a2b0_1sc(din_6_ab0_1sc), .a2b1_1sc(din_6_ab1_1sc),
           .msk_a2b0(din_6_msk_ab0), .msk_a2b1(din_6_msk_ab1),
           .msk_a2b0_1sc(din_6_msk_ab0_1sc), .msk_a2b1_1sc(din_6_msk_ab1_1sc),
           
           .a3b0(din_8_ab0),
           .a3b0_1sc(din_8_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_3_calc (
           .clk(clk), .sign(din_signs_reg[3]), 
           .p(addr_5_3),
           .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
           .a0b0_1sc(din_3_ab0_1sc), .a0b1_1sc(din_3_ab1_1sc), .a0b2_1sc(din_3_ab2_1sc), .a0b3_1sc(din_3_ab3_1sc),
           .msk_a0b0(din_3_msk_ab0), .msk_a0b1(din_3_msk_ab1), .msk_a0b2(din_3_msk_ab2), .msk_a0b3(din_3_msk_ab3),
           .msk_a0b0_1sc(din_3_msk_ab0_1sc), .msk_a0b1_1sc(din_3_msk_ab1_1sc), .msk_a0b2_1sc(din_3_msk_ab2_1sc), .msk_a0b3_1sc(din_3_msk_ab3_1sc),

           .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2),
           .a1b0_1sc(din_5_ab0_1sc), .a1b1_1sc(din_5_ab1_1sc), .a1b2_1sc(din_5_ab2_1sc),
           .msk_a1b0(din_5_msk_ab0), .msk_a1b1(din_5_msk_ab1), .msk_a1b2(din_5_msk_ab2),
           .msk_a1b0_1sc(din_5_msk_ab0_1sc), .msk_a1b1_1sc(din_5_msk_ab1_1sc), .msk_a1b2_1sc(din_5_msk_ab2_1sc),

           .a2b0(din_7_ab0), .a2b1(din_7_ab1),
           .a2b0_1sc(din_7_ab0_1sc), .a2b1_1sc(din_7_ab1_1sc),
           .msk_a2b0(din_7_msk_ab0), .msk_a2b1(din_7_msk_ab1),
           .msk_a2b0_1sc(din_7_msk_ab0_1sc), .msk_a2b1_1sc(din_7_msk_ab1_1sc),
           
           .a3b0(din_9_ab0),
           .a3b0_1sc(din_9_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_4_calc (
           .clk(clk), .sign(din_signs_reg[4]), 
           .p(addr_5_4),
           .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
           .a0b0_1sc(din_4_ab0_1sc), .a0b1_1sc(din_4_ab1_1sc), .a0b2_1sc(din_4_ab2_1sc), .a0b3_1sc(din_4_ab3_1sc),
           .msk_a0b0(din_4_msk_ab0), .msk_a0b1(din_4_msk_ab1), .msk_a0b2(din_4_msk_ab2), .msk_a0b3(din_4_msk_ab3),
           .msk_a0b0_1sc(din_4_msk_ab0_1sc), .msk_a0b1_1sc(din_4_msk_ab1_1sc), .msk_a0b2_1sc(din_4_msk_ab2_1sc), .msk_a0b3_1sc(din_4_msk_ab3_1sc),

           .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2),
           .a1b0_1sc(din_6_ab0_1sc), .a1b1_1sc(din_6_ab1_1sc), .a1b2_1sc(din_6_ab2_1sc),
           .msk_a1b0(din_6_msk_ab0), .msk_a1b1(din_6_msk_ab1), .msk_a1b2(din_6_msk_ab2),
           .msk_a1b0_1sc(din_6_msk_ab0_1sc), .msk_a1b1_1sc(din_6_msk_ab1_1sc), .msk_a1b2_1sc(din_6_msk_ab2_1sc),

           .a2b0(din_8_ab0), .a2b1(din_8_ab1),
           .a2b0_1sc(din_8_ab0_1sc), .a2b1_1sc(din_8_ab1_1sc),
           .msk_a2b0(din_8_msk_ab0), .msk_a2b1(din_8_msk_ab1),
           .msk_a2b0_1sc(din_8_msk_ab0_1sc), .msk_a2b1_1sc(din_8_msk_ab1_1sc),
           
           .a3b0(din_10_ab0),
           .a3b0_1sc(din_10_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_5_calc (
           .clk(clk), .sign(din_signs_reg[5]), 
           .p(addr_5_5),
           .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
           .a0b0_1sc(din_5_ab0_1sc), .a0b1_1sc(din_5_ab1_1sc), .a0b2_1sc(din_5_ab2_1sc), .a0b3_1sc(din_5_ab3_1sc),
           .msk_a0b0(din_5_msk_ab0), .msk_a0b1(din_5_msk_ab1), .msk_a0b2(din_5_msk_ab2), .msk_a0b3(din_5_msk_ab3),
           .msk_a0b0_1sc(din_5_msk_ab0_1sc), .msk_a0b1_1sc(din_5_msk_ab1_1sc), .msk_a0b2_1sc(din_5_msk_ab2_1sc), .msk_a0b3_1sc(din_5_msk_ab3_1sc),

           .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2),
           .a1b0_1sc(din_7_ab0_1sc), .a1b1_1sc(din_7_ab1_1sc), .a1b2_1sc(din_7_ab2_1sc),
           .msk_a1b0(din_7_msk_ab0), .msk_a1b1(din_7_msk_ab1), .msk_a1b2(din_7_msk_ab2),
           .msk_a1b0_1sc(din_7_msk_ab0_1sc), .msk_a1b1_1sc(din_7_msk_ab1_1sc), .msk_a1b2_1sc(din_7_msk_ab2_1sc),

           .a2b0(din_9_ab0), .a2b1(din_9_ab1),
           .a2b0_1sc(din_9_ab0_1sc), .a2b1_1sc(din_9_ab1_1sc),
           .msk_a2b0(din_9_msk_ab0), .msk_a2b1(din_9_msk_ab1),
           .msk_a2b0_1sc(din_9_msk_ab0_1sc), .msk_a2b1_1sc(din_9_msk_ab1_1sc),
           
           .a3b0(din_11_ab0),
           .a3b0_1sc(din_11_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_6_calc (
           .clk(clk), .sign(din_signs_reg[6]), 
           .p(addr_5_6),
           .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
           .a0b0_1sc(din_6_ab0_1sc), .a0b1_1sc(din_6_ab1_1sc), .a0b2_1sc(din_6_ab2_1sc), .a0b3_1sc(din_6_ab3_1sc),
           .msk_a0b0(din_6_msk_ab0), .msk_a0b1(din_6_msk_ab1), .msk_a0b2(din_6_msk_ab2), .msk_a0b3(din_6_msk_ab3),
           .msk_a0b0_1sc(din_6_msk_ab0_1sc), .msk_a0b1_1sc(din_6_msk_ab1_1sc), .msk_a0b2_1sc(din_6_msk_ab2_1sc), .msk_a0b3_1sc(din_6_msk_ab3_1sc),

           .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2),
           .a1b0_1sc(din_8_ab0_1sc), .a1b1_1sc(din_8_ab1_1sc), .a1b2_1sc(din_8_ab2_1sc),
           .msk_a1b0(din_8_msk_ab0), .msk_a1b1(din_8_msk_ab1), .msk_a1b2(din_8_msk_ab2),
           .msk_a1b0_1sc(din_8_msk_ab0_1sc), .msk_a1b1_1sc(din_8_msk_ab1_1sc), .msk_a1b2_1sc(din_8_msk_ab2_1sc),

           .a2b0(din_10_ab0), .a2b1(din_10_ab1),
           .a2b0_1sc(din_10_ab0_1sc), .a2b1_1sc(din_10_ab1_1sc),
           .msk_a2b0(din_10_msk_ab0), .msk_a2b1(din_10_msk_ab1),
           .msk_a2b0_1sc(din_10_msk_ab0_1sc), .msk_a2b1_1sc(din_10_msk_ab1_1sc),
           
           .a3b0(din_12_ab0),
           .a3b0_1sc(din_12_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_7_calc (
           .clk(clk), .sign(din_signs_reg[7]), 
           .p(addr_5_7),
           .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
           .a0b0_1sc(din_7_ab0_1sc), .a0b1_1sc(din_7_ab1_1sc), .a0b2_1sc(din_7_ab2_1sc), .a0b3_1sc(din_7_ab3_1sc),
           .msk_a0b0(din_7_msk_ab0), .msk_a0b1(din_7_msk_ab1), .msk_a0b2(din_7_msk_ab2), .msk_a0b3(din_7_msk_ab3),
           .msk_a0b0_1sc(din_7_msk_ab0_1sc), .msk_a0b1_1sc(din_7_msk_ab1_1sc), .msk_a0b2_1sc(din_7_msk_ab2_1sc), .msk_a0b3_1sc(din_7_msk_ab3_1sc),

           .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2),
           .a1b0_1sc(din_9_ab0_1sc), .a1b1_1sc(din_9_ab1_1sc), .a1b2_1sc(din_9_ab2_1sc),
           .msk_a1b0(din_9_msk_ab0), .msk_a1b1(din_9_msk_ab1), .msk_a1b2(din_9_msk_ab2),
           .msk_a1b0_1sc(din_9_msk_ab0_1sc), .msk_a1b1_1sc(din_9_msk_ab1_1sc), .msk_a1b2_1sc(din_9_msk_ab2_1sc),

           .a2b0(din_11_ab0), .a2b1(din_11_ab1),
           .a2b0_1sc(din_11_ab0_1sc), .a2b1_1sc(din_11_ab1_1sc),
           .msk_a2b0(din_11_msk_ab0), .msk_a2b1(din_11_msk_ab1),
           .msk_a2b0_1sc(din_11_msk_ab0_1sc), .msk_a2b1_1sc(din_11_msk_ab1_1sc),
           
           .a3b0(din_13_ab0),
           .a3b0_1sc(din_13_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_8_calc (
           .clk(clk), .sign(din_signs_reg[8]), 
           .p(addr_5_8),
           .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
           .a0b0_1sc(din_8_ab0_1sc), .a0b1_1sc(din_8_ab1_1sc), .a0b2_1sc(din_8_ab2_1sc), .a0b3_1sc(din_8_ab3_1sc),
           .msk_a0b0(din_8_msk_ab0), .msk_a0b1(din_8_msk_ab1), .msk_a0b2(din_8_msk_ab2), .msk_a0b3(din_8_msk_ab3),
           .msk_a0b0_1sc(din_8_msk_ab0_1sc), .msk_a0b1_1sc(din_8_msk_ab1_1sc), .msk_a0b2_1sc(din_8_msk_ab2_1sc), .msk_a0b3_1sc(din_8_msk_ab3_1sc),

           .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2),
           .a1b0_1sc(din_10_ab0_1sc), .a1b1_1sc(din_10_ab1_1sc), .a1b2_1sc(din_10_ab2_1sc),
           .msk_a1b0(din_10_msk_ab0), .msk_a1b1(din_10_msk_ab1), .msk_a1b2(din_10_msk_ab2),
           .msk_a1b0_1sc(din_10_msk_ab0_1sc), .msk_a1b1_1sc(din_10_msk_ab1_1sc), .msk_a1b2_1sc(din_10_msk_ab2_1sc),

           .a2b0(din_12_ab0), .a2b1(din_12_ab1),
           .a2b0_1sc(din_12_ab0_1sc), .a2b1_1sc(din_12_ab1_1sc),
           .msk_a2b0(din_12_msk_ab0), .msk_a2b1(din_12_msk_ab1),
           .msk_a2b0_1sc(din_12_msk_ab0_1sc), .msk_a2b1_1sc(din_12_msk_ab1_1sc),
           
           .a3b0(din_14_ab0),
           .a3b0_1sc(din_14_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_9_calc (
           .clk(clk), .sign(din_signs_reg[9]), 
           .p(addr_5_9),
           .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
           .a0b0_1sc(din_9_ab0_1sc), .a0b1_1sc(din_9_ab1_1sc), .a0b2_1sc(din_9_ab2_1sc), .a0b3_1sc(din_9_ab3_1sc),
           .msk_a0b0(din_9_msk_ab0), .msk_a0b1(din_9_msk_ab1), .msk_a0b2(din_9_msk_ab2), .msk_a0b3(din_9_msk_ab3),
           .msk_a0b0_1sc(din_9_msk_ab0_1sc), .msk_a0b1_1sc(din_9_msk_ab1_1sc), .msk_a0b2_1sc(din_9_msk_ab2_1sc), .msk_a0b3_1sc(din_9_msk_ab3_1sc),

           .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2),
           .a1b0_1sc(din_11_ab0_1sc), .a1b1_1sc(din_11_ab1_1sc), .a1b2_1sc(din_11_ab2_1sc),
           .msk_a1b0(din_11_msk_ab0), .msk_a1b1(din_11_msk_ab1), .msk_a1b2(din_11_msk_ab2),
           .msk_a1b0_1sc(din_11_msk_ab0_1sc), .msk_a1b1_1sc(din_11_msk_ab1_1sc), .msk_a1b2_1sc(din_11_msk_ab2_1sc),

           .a2b0(din_13_ab0), .a2b1(din_13_ab1),
           .a2b0_1sc(din_13_ab0_1sc), .a2b1_1sc(din_13_ab1_1sc),
           .msk_a2b0(din_13_msk_ab0), .msk_a2b1(din_13_msk_ab1),
           .msk_a2b0_1sc(din_13_msk_ab0_1sc), .msk_a2b1_1sc(din_13_msk_ab1_1sc),
           
           .a3b0(din_15_ab0),
           .a3b0_1sc(din_15_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_10_calc (
           .clk(clk), .sign(din_signs_reg[10]), 
           .p(addr_5_10),
           .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
           .a0b0_1sc(din_10_ab0_1sc), .a0b1_1sc(din_10_ab1_1sc), .a0b2_1sc(din_10_ab2_1sc), .a0b3_1sc(din_10_ab3_1sc),
           .msk_a0b0(din_10_msk_ab0), .msk_a0b1(din_10_msk_ab1), .msk_a0b2(din_10_msk_ab2), .msk_a0b3(din_10_msk_ab3),
           .msk_a0b0_1sc(din_10_msk_ab0_1sc), .msk_a0b1_1sc(din_10_msk_ab1_1sc), .msk_a0b2_1sc(din_10_msk_ab2_1sc), .msk_a0b3_1sc(din_10_msk_ab3_1sc),

           .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2),
           .a1b0_1sc(din_12_ab0_1sc), .a1b1_1sc(din_12_ab1_1sc), .a1b2_1sc(din_12_ab2_1sc),
           .msk_a1b0(din_12_msk_ab0), .msk_a1b1(din_12_msk_ab1), .msk_a1b2(din_12_msk_ab2),
           .msk_a1b0_1sc(din_12_msk_ab0_1sc), .msk_a1b1_1sc(din_12_msk_ab1_1sc), .msk_a1b2_1sc(din_12_msk_ab2_1sc),

           .a2b0(din_14_ab0), .a2b1(din_14_ab1),
           .a2b0_1sc(din_14_ab0_1sc), .a2b1_1sc(din_14_ab1_1sc),
           .msk_a2b0(din_14_msk_ab0), .msk_a2b1(din_14_msk_ab1),
           .msk_a2b0_1sc(din_14_msk_ab0_1sc), .msk_a2b1_1sc(din_14_msk_ab1_1sc),
           
           .a3b0(din_16_ab0),
           .a3b0_1sc(din_16_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_11_calc (
           .clk(clk), .sign(din_signs_reg[11]), 
           .p(addr_5_11),
           .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
           .a0b0_1sc(din_11_ab0_1sc), .a0b1_1sc(din_11_ab1_1sc), .a0b2_1sc(din_11_ab2_1sc), .a0b3_1sc(din_11_ab3_1sc),
           .msk_a0b0(din_11_msk_ab0), .msk_a0b1(din_11_msk_ab1), .msk_a0b2(din_11_msk_ab2), .msk_a0b3(din_11_msk_ab3),
           .msk_a0b0_1sc(din_11_msk_ab0_1sc), .msk_a0b1_1sc(din_11_msk_ab1_1sc), .msk_a0b2_1sc(din_11_msk_ab2_1sc), .msk_a0b3_1sc(din_11_msk_ab3_1sc),

           .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2),
           .a1b0_1sc(din_13_ab0_1sc), .a1b1_1sc(din_13_ab1_1sc), .a1b2_1sc(din_13_ab2_1sc),
           .msk_a1b0(din_13_msk_ab0), .msk_a1b1(din_13_msk_ab1), .msk_a1b2(din_13_msk_ab2),
           .msk_a1b0_1sc(din_13_msk_ab0_1sc), .msk_a1b1_1sc(din_13_msk_ab1_1sc), .msk_a1b2_1sc(din_13_msk_ab2_1sc),

           .a2b0(din_15_ab0), .a2b1(din_15_ab1),
           .a2b0_1sc(din_15_ab0_1sc), .a2b1_1sc(din_15_ab1_1sc),
           .msk_a2b0(din_15_msk_ab0), .msk_a2b1(din_15_msk_ab1),
           .msk_a2b0_1sc(din_15_msk_ab0_1sc), .msk_a2b1_1sc(din_15_msk_ab1_1sc),
           
           .a3b0(din_17_ab0),
           .a3b0_1sc(din_17_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_12_calc (
           .clk(clk), .sign(din_signs_reg[12]), 
           .p(addr_5_12),
           .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
           .a0b0_1sc(din_12_ab0_1sc), .a0b1_1sc(din_12_ab1_1sc), .a0b2_1sc(din_12_ab2_1sc), .a0b3_1sc(din_12_ab3_1sc),
           .msk_a0b0(din_12_msk_ab0), .msk_a0b1(din_12_msk_ab1), .msk_a0b2(din_12_msk_ab2), .msk_a0b3(din_12_msk_ab3),
           .msk_a0b0_1sc(din_12_msk_ab0_1sc), .msk_a0b1_1sc(din_12_msk_ab1_1sc), .msk_a0b2_1sc(din_12_msk_ab2_1sc), .msk_a0b3_1sc(din_12_msk_ab3_1sc),

           .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2),
           .a1b0_1sc(din_14_ab0_1sc), .a1b1_1sc(din_14_ab1_1sc), .a1b2_1sc(din_14_ab2_1sc),
           .msk_a1b0(din_14_msk_ab0), .msk_a1b1(din_14_msk_ab1), .msk_a1b2(din_14_msk_ab2),
           .msk_a1b0_1sc(din_14_msk_ab0_1sc), .msk_a1b1_1sc(din_14_msk_ab1_1sc), .msk_a1b2_1sc(din_14_msk_ab2_1sc),

           .a2b0(din_16_ab0), .a2b1(din_16_ab1),
           .a2b0_1sc(din_16_ab0_1sc), .a2b1_1sc(din_16_ab1_1sc),
           .msk_a2b0(din_16_msk_ab0), .msk_a2b1(din_16_msk_ab1),
           .msk_a2b0_1sc(din_16_msk_ab0_1sc), .msk_a2b1_1sc(din_16_msk_ab1_1sc),
           
           .a3b0(din_18_ab0),
           .a3b0_1sc(din_18_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_13_calc (
           .clk(clk), .sign(din_signs_reg[13]), 
           .p(addr_5_13),
           .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
           .a0b0_1sc(din_13_ab0_1sc), .a0b1_1sc(din_13_ab1_1sc), .a0b2_1sc(din_13_ab2_1sc), .a0b3_1sc(din_13_ab3_1sc),
           .msk_a0b0(din_13_msk_ab0), .msk_a0b1(din_13_msk_ab1), .msk_a0b2(din_13_msk_ab2), .msk_a0b3(din_13_msk_ab3),
           .msk_a0b0_1sc(din_13_msk_ab0_1sc), .msk_a0b1_1sc(din_13_msk_ab1_1sc), .msk_a0b2_1sc(din_13_msk_ab2_1sc), .msk_a0b3_1sc(din_13_msk_ab3_1sc),

           .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2),
           .a1b0_1sc(din_15_ab0_1sc), .a1b1_1sc(din_15_ab1_1sc), .a1b2_1sc(din_15_ab2_1sc),
           .msk_a1b0(din_15_msk_ab0), .msk_a1b1(din_15_msk_ab1), .msk_a1b2(din_15_msk_ab2),
           .msk_a1b0_1sc(din_15_msk_ab0_1sc), .msk_a1b1_1sc(din_15_msk_ab1_1sc), .msk_a1b2_1sc(din_15_msk_ab2_1sc),

           .a2b0(din_17_ab0), .a2b1(din_17_ab1),
           .a2b0_1sc(din_17_ab0_1sc), .a2b1_1sc(din_17_ab1_1sc),
           .msk_a2b0(din_17_msk_ab0), .msk_a2b1(din_17_msk_ab1),
           .msk_a2b0_1sc(din_17_msk_ab0_1sc), .msk_a2b1_1sc(din_17_msk_ab1_1sc),
           
           .a3b0(din_19_ab0),
           .a3b0_1sc(din_19_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_14_calc (
           .clk(clk), .sign(din_signs_reg[14]), 
           .p(addr_5_14),
           .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
           .a0b0_1sc(din_14_ab0_1sc), .a0b1_1sc(din_14_ab1_1sc), .a0b2_1sc(din_14_ab2_1sc), .a0b3_1sc(din_14_ab3_1sc),
           .msk_a0b0(din_14_msk_ab0), .msk_a0b1(din_14_msk_ab1), .msk_a0b2(din_14_msk_ab2), .msk_a0b3(din_14_msk_ab3),
           .msk_a0b0_1sc(din_14_msk_ab0_1sc), .msk_a0b1_1sc(din_14_msk_ab1_1sc), .msk_a0b2_1sc(din_14_msk_ab2_1sc), .msk_a0b3_1sc(din_14_msk_ab3_1sc),

           .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2),
           .a1b0_1sc(din_16_ab0_1sc), .a1b1_1sc(din_16_ab1_1sc), .a1b2_1sc(din_16_ab2_1sc),
           .msk_a1b0(din_16_msk_ab0), .msk_a1b1(din_16_msk_ab1), .msk_a1b2(din_16_msk_ab2),
           .msk_a1b0_1sc(din_16_msk_ab0_1sc), .msk_a1b1_1sc(din_16_msk_ab1_1sc), .msk_a1b2_1sc(din_16_msk_ab2_1sc),

           .a2b0(din_18_ab0), .a2b1(din_18_ab1),
           .a2b0_1sc(din_18_ab0_1sc), .a2b1_1sc(din_18_ab1_1sc),
           .msk_a2b0(din_18_msk_ab0), .msk_a2b1(din_18_msk_ab1),
           .msk_a2b0_1sc(din_18_msk_ab0_1sc), .msk_a2b1_1sc(din_18_msk_ab1_1sc),
           
           .a3b0(din_20_ab0),
           .a3b0_1sc(din_20_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_15_calc (
           .clk(clk), .sign(din_signs_reg[15]), 
           .p(addr_5_15),
           .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
           .a0b0_1sc(din_15_ab0_1sc), .a0b1_1sc(din_15_ab1_1sc), .a0b2_1sc(din_15_ab2_1sc), .a0b3_1sc(din_15_ab3_1sc),
           .msk_a0b0(din_15_msk_ab0), .msk_a0b1(din_15_msk_ab1), .msk_a0b2(din_15_msk_ab2), .msk_a0b3(din_15_msk_ab3),
           .msk_a0b0_1sc(din_15_msk_ab0_1sc), .msk_a0b1_1sc(din_15_msk_ab1_1sc), .msk_a0b2_1sc(din_15_msk_ab2_1sc), .msk_a0b3_1sc(din_15_msk_ab3_1sc),

           .a1b0(din_17_ab0), .a1b1(din_17_ab1), .a1b2(din_17_ab2),
           .a1b0_1sc(din_17_ab0_1sc), .a1b1_1sc(din_17_ab1_1sc), .a1b2_1sc(din_17_ab2_1sc),
           .msk_a1b0(din_17_msk_ab0), .msk_a1b1(din_17_msk_ab1), .msk_a1b2(din_17_msk_ab2),
           .msk_a1b0_1sc(din_17_msk_ab0_1sc), .msk_a1b1_1sc(din_17_msk_ab1_1sc), .msk_a1b2_1sc(din_17_msk_ab2_1sc),

           .a2b0(din_19_ab0), .a2b1(din_19_ab1),
           .a2b0_1sc(din_19_ab0_1sc), .a2b1_1sc(din_19_ab1_1sc),
           .msk_a2b0(din_19_msk_ab0), .msk_a2b1(din_19_msk_ab1),
           .msk_a2b0_1sc(din_19_msk_ab0_1sc), .msk_a2b1_1sc(din_19_msk_ab1_1sc),
           
           .a3b0(din_21_ab0),
           .a3b0_1sc(din_21_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_16_calc (
           .clk(clk), .sign(din_signs_reg[16]), 
           .p(addr_5_16),
           .a0b0(din_16_ab0), .a0b1(din_16_ab1), .a0b2(din_16_ab2), .a0b3(din_16_ab3),
           .a0b0_1sc(din_16_ab0_1sc), .a0b1_1sc(din_16_ab1_1sc), .a0b2_1sc(din_16_ab2_1sc), .a0b3_1sc(din_16_ab3_1sc),
           .msk_a0b0(din_16_msk_ab0), .msk_a0b1(din_16_msk_ab1), .msk_a0b2(din_16_msk_ab2), .msk_a0b3(din_16_msk_ab3),
           .msk_a0b0_1sc(din_16_msk_ab0_1sc), .msk_a0b1_1sc(din_16_msk_ab1_1sc), .msk_a0b2_1sc(din_16_msk_ab2_1sc), .msk_a0b3_1sc(din_16_msk_ab3_1sc),

           .a1b0(din_18_ab0), .a1b1(din_18_ab1), .a1b2(din_18_ab2),
           .a1b0_1sc(din_18_ab0_1sc), .a1b1_1sc(din_18_ab1_1sc), .a1b2_1sc(din_18_ab2_1sc),
           .msk_a1b0(din_18_msk_ab0), .msk_a1b1(din_18_msk_ab1), .msk_a1b2(din_18_msk_ab2),
           .msk_a1b0_1sc(din_18_msk_ab0_1sc), .msk_a1b1_1sc(din_18_msk_ab1_1sc), .msk_a1b2_1sc(din_18_msk_ab2_1sc),

           .a2b0(din_20_ab0), .a2b1(din_20_ab1),
           .a2b0_1sc(din_20_ab0_1sc), .a2b1_1sc(din_20_ab1_1sc),
           .msk_a2b0(din_20_msk_ab0), .msk_a2b1(din_20_msk_ab1),
           .msk_a2b0_1sc(din_20_msk_ab0_1sc), .msk_a2b1_1sc(din_20_msk_ab1_1sc),
           
           .a3b0(din_22_ab0),
           .a3b0_1sc(din_22_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_17_calc (
           .clk(clk), .sign(din_signs_reg[17]), 
           .p(addr_5_17),
           .a0b0(din_17_ab0), .a0b1(din_17_ab1), .a0b2(din_17_ab2), .a0b3(din_17_ab3),
           .a0b0_1sc(din_17_ab0_1sc), .a0b1_1sc(din_17_ab1_1sc), .a0b2_1sc(din_17_ab2_1sc), .a0b3_1sc(din_17_ab3_1sc),
           .msk_a0b0(din_17_msk_ab0), .msk_a0b1(din_17_msk_ab1), .msk_a0b2(din_17_msk_ab2), .msk_a0b3(din_17_msk_ab3),
           .msk_a0b0_1sc(din_17_msk_ab0_1sc), .msk_a0b1_1sc(din_17_msk_ab1_1sc), .msk_a0b2_1sc(din_17_msk_ab2_1sc), .msk_a0b3_1sc(din_17_msk_ab3_1sc),

           .a1b0(din_19_ab0), .a1b1(din_19_ab1), .a1b2(din_19_ab2),
           .a1b0_1sc(din_19_ab0_1sc), .a1b1_1sc(din_19_ab1_1sc), .a1b2_1sc(din_19_ab2_1sc),
           .msk_a1b0(din_19_msk_ab0), .msk_a1b1(din_19_msk_ab1), .msk_a1b2(din_19_msk_ab2),
           .msk_a1b0_1sc(din_19_msk_ab0_1sc), .msk_a1b1_1sc(din_19_msk_ab1_1sc), .msk_a1b2_1sc(din_19_msk_ab2_1sc),

           .a2b0(din_21_ab0), .a2b1(din_21_ab1),
           .a2b0_1sc(din_21_ab0_1sc), .a2b1_1sc(din_21_ab1_1sc),
           .msk_a2b0(din_21_msk_ab0), .msk_a2b1(din_21_msk_ab1),
           .msk_a2b0_1sc(din_21_msk_ab0_1sc), .msk_a2b1_1sc(din_21_msk_ab1_1sc),
           
           .a3b0(din_23_ab0),
           .a3b0_1sc(din_23_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_18_calc (
           .clk(clk), .sign(din_signs_reg[18]), 
           .p(addr_5_18),
           .a0b0(din_18_ab0), .a0b1(din_18_ab1), .a0b2(din_18_ab2), .a0b3(din_18_ab3),
           .a0b0_1sc(din_18_ab0_1sc), .a0b1_1sc(din_18_ab1_1sc), .a0b2_1sc(din_18_ab2_1sc), .a0b3_1sc(din_18_ab3_1sc),
           .msk_a0b0(din_18_msk_ab0), .msk_a0b1(din_18_msk_ab1), .msk_a0b2(din_18_msk_ab2), .msk_a0b3(din_18_msk_ab3),
           .msk_a0b0_1sc(din_18_msk_ab0_1sc), .msk_a0b1_1sc(din_18_msk_ab1_1sc), .msk_a0b2_1sc(din_18_msk_ab2_1sc), .msk_a0b3_1sc(din_18_msk_ab3_1sc),

           .a1b0(din_20_ab0), .a1b1(din_20_ab1), .a1b2(din_20_ab2),
           .a1b0_1sc(din_20_ab0_1sc), .a1b1_1sc(din_20_ab1_1sc), .a1b2_1sc(din_20_ab2_1sc),
           .msk_a1b0(din_20_msk_ab0), .msk_a1b1(din_20_msk_ab1), .msk_a1b2(din_20_msk_ab2),
           .msk_a1b0_1sc(din_20_msk_ab0_1sc), .msk_a1b1_1sc(din_20_msk_ab1_1sc), .msk_a1b2_1sc(din_20_msk_ab2_1sc),

           .a2b0(din_22_ab0), .a2b1(din_22_ab1),
           .a2b0_1sc(din_22_ab0_1sc), .a2b1_1sc(din_22_ab1_1sc),
           .msk_a2b0(din_22_msk_ab0), .msk_a2b1(din_22_msk_ab1),
           .msk_a2b0_1sc(din_22_msk_ab0_1sc), .msk_a2b1_1sc(din_22_msk_ab1_1sc),
           
           .a3b0(din_24_ab0),
           .a3b0_1sc(din_24_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_19_calc (
           .clk(clk), .sign(din_signs_reg[19]), 
           .p(addr_5_19),
           .a0b0(din_19_ab0), .a0b1(din_19_ab1), .a0b2(din_19_ab2), .a0b3(din_19_ab3),
           .a0b0_1sc(din_19_ab0_1sc), .a0b1_1sc(din_19_ab1_1sc), .a0b2_1sc(din_19_ab2_1sc), .a0b3_1sc(din_19_ab3_1sc),
           .msk_a0b0(din_19_msk_ab0), .msk_a0b1(din_19_msk_ab1), .msk_a0b2(din_19_msk_ab2), .msk_a0b3(din_19_msk_ab3),
           .msk_a0b0_1sc(din_19_msk_ab0_1sc), .msk_a0b1_1sc(din_19_msk_ab1_1sc), .msk_a0b2_1sc(din_19_msk_ab2_1sc), .msk_a0b3_1sc(din_19_msk_ab3_1sc),

           .a1b0(din_21_ab0), .a1b1(din_21_ab1), .a1b2(din_21_ab2),
           .a1b0_1sc(din_21_ab0_1sc), .a1b1_1sc(din_21_ab1_1sc), .a1b2_1sc(din_21_ab2_1sc),
           .msk_a1b0(din_21_msk_ab0), .msk_a1b1(din_21_msk_ab1), .msk_a1b2(din_21_msk_ab2),
           .msk_a1b0_1sc(din_21_msk_ab0_1sc), .msk_a1b1_1sc(din_21_msk_ab1_1sc), .msk_a1b2_1sc(din_21_msk_ab2_1sc),

           .a2b0(din_23_ab0), .a2b1(din_23_ab1),
           .a2b0_1sc(din_23_ab0_1sc), .a2b1_1sc(din_23_ab1_1sc),
           .msk_a2b0(din_23_msk_ab0), .msk_a2b1(din_23_msk_ab1),
           .msk_a2b0_1sc(din_23_msk_ab0_1sc), .msk_a2b1_1sc(din_23_msk_ab1_1sc),
           
           .a3b0(din_25_ab0),
           .a3b0_1sc(din_25_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_20_calc (
           .clk(clk), .sign(din_signs_reg[20]), 
           .p(addr_5_20),
           .a0b0(din_20_ab0), .a0b1(din_20_ab1), .a0b2(din_20_ab2), .a0b3(din_20_ab3),
           .a0b0_1sc(din_20_ab0_1sc), .a0b1_1sc(din_20_ab1_1sc), .a0b2_1sc(din_20_ab2_1sc), .a0b3_1sc(din_20_ab3_1sc),
           .msk_a0b0(din_20_msk_ab0), .msk_a0b1(din_20_msk_ab1), .msk_a0b2(din_20_msk_ab2), .msk_a0b3(din_20_msk_ab3),
           .msk_a0b0_1sc(din_20_msk_ab0_1sc), .msk_a0b1_1sc(din_20_msk_ab1_1sc), .msk_a0b2_1sc(din_20_msk_ab2_1sc), .msk_a0b3_1sc(din_20_msk_ab3_1sc),

           .a1b0(din_22_ab0), .a1b1(din_22_ab1), .a1b2(din_22_ab2),
           .a1b0_1sc(din_22_ab0_1sc), .a1b1_1sc(din_22_ab1_1sc), .a1b2_1sc(din_22_ab2_1sc),
           .msk_a1b0(din_22_msk_ab0), .msk_a1b1(din_22_msk_ab1), .msk_a1b2(din_22_msk_ab2),
           .msk_a1b0_1sc(din_22_msk_ab0_1sc), .msk_a1b1_1sc(din_22_msk_ab1_1sc), .msk_a1b2_1sc(din_22_msk_ab2_1sc),

           .a2b0(din_24_ab0), .a2b1(din_24_ab1),
           .a2b0_1sc(din_24_ab0_1sc), .a2b1_1sc(din_24_ab1_1sc),
           .msk_a2b0(din_24_msk_ab0), .msk_a2b1(din_24_msk_ab1),
           .msk_a2b0_1sc(din_24_msk_ab0_1sc), .msk_a2b1_1sc(din_24_msk_ab1_1sc),
           
           .a3b0(din_26_ab0),
           .a3b0_1sc(din_26_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_21_calc (
           .clk(clk), .sign(din_signs_reg[21]), 
           .p(addr_5_21),
           .a0b0(din_21_ab0), .a0b1(din_21_ab1), .a0b2(din_21_ab2), .a0b3(din_21_ab3),
           .a0b0_1sc(din_21_ab0_1sc), .a0b1_1sc(din_21_ab1_1sc), .a0b2_1sc(din_21_ab2_1sc), .a0b3_1sc(din_21_ab3_1sc),
           .msk_a0b0(din_21_msk_ab0), .msk_a0b1(din_21_msk_ab1), .msk_a0b2(din_21_msk_ab2), .msk_a0b3(din_21_msk_ab3),
           .msk_a0b0_1sc(din_21_msk_ab0_1sc), .msk_a0b1_1sc(din_21_msk_ab1_1sc), .msk_a0b2_1sc(din_21_msk_ab2_1sc), .msk_a0b3_1sc(din_21_msk_ab3_1sc),

           .a1b0(din_23_ab0), .a1b1(din_23_ab1), .a1b2(din_23_ab2),
           .a1b0_1sc(din_23_ab0_1sc), .a1b1_1sc(din_23_ab1_1sc), .a1b2_1sc(din_23_ab2_1sc),
           .msk_a1b0(din_23_msk_ab0), .msk_a1b1(din_23_msk_ab1), .msk_a1b2(din_23_msk_ab2),
           .msk_a1b0_1sc(din_23_msk_ab0_1sc), .msk_a1b1_1sc(din_23_msk_ab1_1sc), .msk_a1b2_1sc(din_23_msk_ab2_1sc),

           .a2b0(din_25_ab0), .a2b1(din_25_ab1),
           .a2b0_1sc(din_25_ab0_1sc), .a2b1_1sc(din_25_ab1_1sc),
           .msk_a2b0(din_25_msk_ab0), .msk_a2b1(din_25_msk_ab1),
           .msk_a2b0_1sc(din_25_msk_ab0_1sc), .msk_a2b1_1sc(din_25_msk_ab1_1sc),
           
           .a3b0(din_27_ab0),
           .a3b0_1sc(din_27_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_22_calc (
           .clk(clk), .sign(din_signs_reg[22]), 
           .p(addr_5_22),
           .a0b0(din_22_ab0), .a0b1(din_22_ab1), .a0b2(din_22_ab2), .a0b3(din_22_ab3),
           .a0b0_1sc(din_22_ab0_1sc), .a0b1_1sc(din_22_ab1_1sc), .a0b2_1sc(din_22_ab2_1sc), .a0b3_1sc(din_22_ab3_1sc),
           .msk_a0b0(din_22_msk_ab0), .msk_a0b1(din_22_msk_ab1), .msk_a0b2(din_22_msk_ab2), .msk_a0b3(din_22_msk_ab3),
           .msk_a0b0_1sc(din_22_msk_ab0_1sc), .msk_a0b1_1sc(din_22_msk_ab1_1sc), .msk_a0b2_1sc(din_22_msk_ab2_1sc), .msk_a0b3_1sc(din_22_msk_ab3_1sc),

           .a1b0(din_24_ab0), .a1b1(din_24_ab1), .a1b2(din_24_ab2),
           .a1b0_1sc(din_24_ab0_1sc), .a1b1_1sc(din_24_ab1_1sc), .a1b2_1sc(din_24_ab2_1sc),
           .msk_a1b0(din_24_msk_ab0), .msk_a1b1(din_24_msk_ab1), .msk_a1b2(din_24_msk_ab2),
           .msk_a1b0_1sc(din_24_msk_ab0_1sc), .msk_a1b1_1sc(din_24_msk_ab1_1sc), .msk_a1b2_1sc(din_24_msk_ab2_1sc),

           .a2b0(din_26_ab0), .a2b1(din_26_ab1),
           .a2b0_1sc(din_26_ab0_1sc), .a2b1_1sc(din_26_ab1_1sc),
           .msk_a2b0(din_26_msk_ab0), .msk_a2b1(din_26_msk_ab1),
           .msk_a2b0_1sc(din_26_msk_ab0_1sc), .msk_a2b1_1sc(din_26_msk_ab1_1sc),
           
           .a3b0(din_28_ab0),
           .a3b0_1sc(din_28_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_23_calc (
           .clk(clk), .sign(din_signs_reg[23]), 
           .p(addr_5_23),
           .a0b0(din_23_ab0), .a0b1(din_23_ab1), .a0b2(din_23_ab2), .a0b3(din_23_ab3),
           .a0b0_1sc(din_23_ab0_1sc), .a0b1_1sc(din_23_ab1_1sc), .a0b2_1sc(din_23_ab2_1sc), .a0b3_1sc(din_23_ab3_1sc),
           .msk_a0b0(din_23_msk_ab0), .msk_a0b1(din_23_msk_ab1), .msk_a0b2(din_23_msk_ab2), .msk_a0b3(din_23_msk_ab3),
           .msk_a0b0_1sc(din_23_msk_ab0_1sc), .msk_a0b1_1sc(din_23_msk_ab1_1sc), .msk_a0b2_1sc(din_23_msk_ab2_1sc), .msk_a0b3_1sc(din_23_msk_ab3_1sc),

           .a1b0(din_25_ab0), .a1b1(din_25_ab1), .a1b2(din_25_ab2),
           .a1b0_1sc(din_25_ab0_1sc), .a1b1_1sc(din_25_ab1_1sc), .a1b2_1sc(din_25_ab2_1sc),
           .msk_a1b0(din_25_msk_ab0), .msk_a1b1(din_25_msk_ab1), .msk_a1b2(din_25_msk_ab2),
           .msk_a1b0_1sc(din_25_msk_ab0_1sc), .msk_a1b1_1sc(din_25_msk_ab1_1sc), .msk_a1b2_1sc(din_25_msk_ab2_1sc),

           .a2b0(din_27_ab0), .a2b1(din_27_ab1),
           .a2b0_1sc(din_27_ab0_1sc), .a2b1_1sc(din_27_ab1_1sc),
           .msk_a2b0(din_27_msk_ab0), .msk_a2b1(din_27_msk_ab1),
           .msk_a2b0_1sc(din_27_msk_ab0_1sc), .msk_a2b1_1sc(din_27_msk_ab1_1sc),
           
           .a3b0(din_29_ab0),
           .a3b0_1sc(din_29_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_24_calc (
           .clk(clk), .sign(din_signs_reg[24]), 
           .p(addr_5_24),
           .a0b0(din_24_ab0), .a0b1(din_24_ab1), .a0b2(din_24_ab2), .a0b3(din_24_ab3),
           .a0b0_1sc(din_24_ab0_1sc), .a0b1_1sc(din_24_ab1_1sc), .a0b2_1sc(din_24_ab2_1sc), .a0b3_1sc(din_24_ab3_1sc),
           .msk_a0b0(din_24_msk_ab0), .msk_a0b1(din_24_msk_ab1), .msk_a0b2(din_24_msk_ab2), .msk_a0b3(din_24_msk_ab3),
           .msk_a0b0_1sc(din_24_msk_ab0_1sc), .msk_a0b1_1sc(din_24_msk_ab1_1sc), .msk_a0b2_1sc(din_24_msk_ab2_1sc), .msk_a0b3_1sc(din_24_msk_ab3_1sc),

           .a1b0(din_26_ab0), .a1b1(din_26_ab1), .a1b2(din_26_ab2),
           .a1b0_1sc(din_26_ab0_1sc), .a1b1_1sc(din_26_ab1_1sc), .a1b2_1sc(din_26_ab2_1sc),
           .msk_a1b0(din_26_msk_ab0), .msk_a1b1(din_26_msk_ab1), .msk_a1b2(din_26_msk_ab2),
           .msk_a1b0_1sc(din_26_msk_ab0_1sc), .msk_a1b1_1sc(din_26_msk_ab1_1sc), .msk_a1b2_1sc(din_26_msk_ab2_1sc),

           .a2b0(din_28_ab0), .a2b1(din_28_ab1),
           .a2b0_1sc(din_28_ab0_1sc), .a2b1_1sc(din_28_ab1_1sc),
           .msk_a2b0(din_28_msk_ab0), .msk_a2b1(din_28_msk_ab1),
           .msk_a2b0_1sc(din_28_msk_ab0_1sc), .msk_a2b1_1sc(din_28_msk_ab1_1sc),
           
           .a3b0(din_30_ab0),
           .a3b0_1sc(din_30_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_25_calc (
           .clk(clk), .sign(din_signs_reg[25]), 
           .p(addr_5_25),
           .a0b0(din_25_ab0), .a0b1(din_25_ab1), .a0b2(din_25_ab2), .a0b3(din_25_ab3),
           .a0b0_1sc(din_25_ab0_1sc), .a0b1_1sc(din_25_ab1_1sc), .a0b2_1sc(din_25_ab2_1sc), .a0b3_1sc(din_25_ab3_1sc),
           .msk_a0b0(din_25_msk_ab0), .msk_a0b1(din_25_msk_ab1), .msk_a0b2(din_25_msk_ab2), .msk_a0b3(din_25_msk_ab3),
           .msk_a0b0_1sc(din_25_msk_ab0_1sc), .msk_a0b1_1sc(din_25_msk_ab1_1sc), .msk_a0b2_1sc(din_25_msk_ab2_1sc), .msk_a0b3_1sc(din_25_msk_ab3_1sc),

           .a1b0(din_27_ab0), .a1b1(din_27_ab1), .a1b2(din_27_ab2),
           .a1b0_1sc(din_27_ab0_1sc), .a1b1_1sc(din_27_ab1_1sc), .a1b2_1sc(din_27_ab2_1sc),
           .msk_a1b0(din_27_msk_ab0), .msk_a1b1(din_27_msk_ab1), .msk_a1b2(din_27_msk_ab2),
           .msk_a1b0_1sc(din_27_msk_ab0_1sc), .msk_a1b1_1sc(din_27_msk_ab1_1sc), .msk_a1b2_1sc(din_27_msk_ab2_1sc),

           .a2b0(din_29_ab0), .a2b1(din_29_ab1),
           .a2b0_1sc(din_29_ab0_1sc), .a2b1_1sc(din_29_ab1_1sc),
           .msk_a2b0(din_29_msk_ab0), .msk_a2b1(din_29_msk_ab1),
           .msk_a2b0_1sc(din_29_msk_ab0_1sc), .msk_a2b1_1sc(din_29_msk_ab1_1sc),
           
           .a3b0(din_31_ab0),
           .a3b0_1sc(din_31_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_26_calc (
           .clk(clk), .sign(din_signs_reg[26]), 
           .p(addr_5_26),
           .a0b0(din_26_ab0), .a0b1(din_26_ab1), .a0b2(din_26_ab2), .a0b3(din_26_ab3),
           .a0b0_1sc(din_26_ab0_1sc), .a0b1_1sc(din_26_ab1_1sc), .a0b2_1sc(din_26_ab2_1sc), .a0b3_1sc(din_26_ab3_1sc),
           .msk_a0b0(din_26_msk_ab0), .msk_a0b1(din_26_msk_ab1), .msk_a0b2(din_26_msk_ab2), .msk_a0b3(din_26_msk_ab3),
           .msk_a0b0_1sc(din_26_msk_ab0_1sc), .msk_a0b1_1sc(din_26_msk_ab1_1sc), .msk_a0b2_1sc(din_26_msk_ab2_1sc), .msk_a0b3_1sc(din_26_msk_ab3_1sc),

           .a1b0(din_28_ab0), .a1b1(din_28_ab1), .a1b2(din_28_ab2),
           .a1b0_1sc(din_28_ab0_1sc), .a1b1_1sc(din_28_ab1_1sc), .a1b2_1sc(din_28_ab2_1sc),
           .msk_a1b0(din_28_msk_ab0), .msk_a1b1(din_28_msk_ab1), .msk_a1b2(din_28_msk_ab2),
           .msk_a1b0_1sc(din_28_msk_ab0_1sc), .msk_a1b1_1sc(din_28_msk_ab1_1sc), .msk_a1b2_1sc(din_28_msk_ab2_1sc),

           .a2b0(din_30_ab0), .a2b1(din_30_ab1),
           .a2b0_1sc(din_30_ab0_1sc), .a2b1_1sc(din_30_ab1_1sc),
           .msk_a2b0(din_30_msk_ab0), .msk_a2b1(din_30_msk_ab1),
           .msk_a2b0_1sc(din_30_msk_ab0_1sc), .msk_a2b1_1sc(din_30_msk_ab1_1sc),
           
           .a3b0(din_32_ab0),
           .a3b0_1sc(din_32_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_27_calc (
           .clk(clk), .sign(din_signs_reg[27]), 
           .p(addr_5_27),
           .a0b0(din_27_ab0), .a0b1(din_27_ab1), .a0b2(din_27_ab2), .a0b3(din_27_ab3),
           .a0b0_1sc(din_27_ab0_1sc), .a0b1_1sc(din_27_ab1_1sc), .a0b2_1sc(din_27_ab2_1sc), .a0b3_1sc(din_27_ab3_1sc),
           .msk_a0b0(din_27_msk_ab0), .msk_a0b1(din_27_msk_ab1), .msk_a0b2(din_27_msk_ab2), .msk_a0b3(din_27_msk_ab3),
           .msk_a0b0_1sc(din_27_msk_ab0_1sc), .msk_a0b1_1sc(din_27_msk_ab1_1sc), .msk_a0b2_1sc(din_27_msk_ab2_1sc), .msk_a0b3_1sc(din_27_msk_ab3_1sc),

           .a1b0(din_29_ab0), .a1b1(din_29_ab1), .a1b2(din_29_ab2),
           .a1b0_1sc(din_29_ab0_1sc), .a1b1_1sc(din_29_ab1_1sc), .a1b2_1sc(din_29_ab2_1sc),
           .msk_a1b0(din_29_msk_ab0), .msk_a1b1(din_29_msk_ab1), .msk_a1b2(din_29_msk_ab2),
           .msk_a1b0_1sc(din_29_msk_ab0_1sc), .msk_a1b1_1sc(din_29_msk_ab1_1sc), .msk_a1b2_1sc(din_29_msk_ab2_1sc),

           .a2b0(din_31_ab0), .a2b1(din_31_ab1),
           .a2b0_1sc(din_31_ab0_1sc), .a2b1_1sc(din_31_ab1_1sc),
           .msk_a2b0(din_31_msk_ab0), .msk_a2b1(din_31_msk_ab1),
           .msk_a2b0_1sc(din_31_msk_ab0_1sc), .msk_a2b1_1sc(din_31_msk_ab1_1sc),
           
           .a3b0(din_33_ab0),
           .a3b0_1sc(din_33_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_28_calc (
           .clk(clk), .sign(din_signs_reg[28]), 
           .p(addr_5_28),
           .a0b0(din_28_ab0), .a0b1(din_28_ab1), .a0b2(din_28_ab2), .a0b3(din_28_ab3),
           .a0b0_1sc(din_28_ab0_1sc), .a0b1_1sc(din_28_ab1_1sc), .a0b2_1sc(din_28_ab2_1sc), .a0b3_1sc(din_28_ab3_1sc),
           .msk_a0b0(din_28_msk_ab0), .msk_a0b1(din_28_msk_ab1), .msk_a0b2(din_28_msk_ab2), .msk_a0b3(din_28_msk_ab3),
           .msk_a0b0_1sc(din_28_msk_ab0_1sc), .msk_a0b1_1sc(din_28_msk_ab1_1sc), .msk_a0b2_1sc(din_28_msk_ab2_1sc), .msk_a0b3_1sc(din_28_msk_ab3_1sc),

           .a1b0(din_30_ab0), .a1b1(din_30_ab1), .a1b2(din_30_ab2),
           .a1b0_1sc(din_30_ab0_1sc), .a1b1_1sc(din_30_ab1_1sc), .a1b2_1sc(din_30_ab2_1sc),
           .msk_a1b0(din_30_msk_ab0), .msk_a1b1(din_30_msk_ab1), .msk_a1b2(din_30_msk_ab2),
           .msk_a1b0_1sc(din_30_msk_ab0_1sc), .msk_a1b1_1sc(din_30_msk_ab1_1sc), .msk_a1b2_1sc(din_30_msk_ab2_1sc),

           .a2b0(din_32_ab0), .a2b1(din_32_ab1),
           .a2b0_1sc(din_32_ab0_1sc), .a2b1_1sc(din_32_ab1_1sc),
           .msk_a2b0(din_32_msk_ab0), .msk_a2b1(din_32_msk_ab1),
           .msk_a2b0_1sc(din_32_msk_ab0_1sc), .msk_a2b1_1sc(din_32_msk_ab1_1sc),
           
           .a3b0(din_34_ab0),
           .a3b0_1sc(din_34_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_29_calc (
           .clk(clk), .sign(din_signs_reg[29]), 
           .p(addr_5_29),
           .a0b0(din_29_ab0), .a0b1(din_29_ab1), .a0b2(din_29_ab2), .a0b3(din_29_ab3),
           .a0b0_1sc(din_29_ab0_1sc), .a0b1_1sc(din_29_ab1_1sc), .a0b2_1sc(din_29_ab2_1sc), .a0b3_1sc(din_29_ab3_1sc),
           .msk_a0b0(din_29_msk_ab0), .msk_a0b1(din_29_msk_ab1), .msk_a0b2(din_29_msk_ab2), .msk_a0b3(din_29_msk_ab3),
           .msk_a0b0_1sc(din_29_msk_ab0_1sc), .msk_a0b1_1sc(din_29_msk_ab1_1sc), .msk_a0b2_1sc(din_29_msk_ab2_1sc), .msk_a0b3_1sc(din_29_msk_ab3_1sc),

           .a1b0(din_31_ab0), .a1b1(din_31_ab1), .a1b2(din_31_ab2),
           .a1b0_1sc(din_31_ab0_1sc), .a1b1_1sc(din_31_ab1_1sc), .a1b2_1sc(din_31_ab2_1sc),
           .msk_a1b0(din_31_msk_ab0), .msk_a1b1(din_31_msk_ab1), .msk_a1b2(din_31_msk_ab2),
           .msk_a1b0_1sc(din_31_msk_ab0_1sc), .msk_a1b1_1sc(din_31_msk_ab1_1sc), .msk_a1b2_1sc(din_31_msk_ab2_1sc),

           .a2b0(din_33_ab0), .a2b1(din_33_ab1),
           .a2b0_1sc(din_33_ab0_1sc), .a2b1_1sc(din_33_ab1_1sc),
           .msk_a2b0(din_33_msk_ab0), .msk_a2b1(din_33_msk_ab1),
           .msk_a2b0_1sc(din_33_msk_ab0_1sc), .msk_a2b1_1sc(din_33_msk_ab1_1sc),
           
           .a3b0(din_35_ab0),
           .a3b0_1sc(din_35_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_30_calc (
           .clk(clk), .sign(din_signs_reg[30]), 
           .p(addr_5_30),
           .a0b0(din_30_ab0), .a0b1(din_30_ab1), .a0b2(din_30_ab2), .a0b3(din_30_ab3),
           .a0b0_1sc(din_30_ab0_1sc), .a0b1_1sc(din_30_ab1_1sc), .a0b2_1sc(din_30_ab2_1sc), .a0b3_1sc(din_30_ab3_1sc),
           .msk_a0b0(din_30_msk_ab0), .msk_a0b1(din_30_msk_ab1), .msk_a0b2(din_30_msk_ab2), .msk_a0b3(din_30_msk_ab3),
           .msk_a0b0_1sc(din_30_msk_ab0_1sc), .msk_a0b1_1sc(din_30_msk_ab1_1sc), .msk_a0b2_1sc(din_30_msk_ab2_1sc), .msk_a0b3_1sc(din_30_msk_ab3_1sc),

           .a1b0(din_32_ab0), .a1b1(din_32_ab1), .a1b2(din_32_ab2),
           .a1b0_1sc(din_32_ab0_1sc), .a1b1_1sc(din_32_ab1_1sc), .a1b2_1sc(din_32_ab2_1sc),
           .msk_a1b0(din_32_msk_ab0), .msk_a1b1(din_32_msk_ab1), .msk_a1b2(din_32_msk_ab2),
           .msk_a1b0_1sc(din_32_msk_ab0_1sc), .msk_a1b1_1sc(din_32_msk_ab1_1sc), .msk_a1b2_1sc(din_32_msk_ab2_1sc),

           .a2b0(din_34_ab0), .a2b1(din_34_ab1),
           .a2b0_1sc(din_34_ab0_1sc), .a2b1_1sc(din_34_ab1_1sc),
           .msk_a2b0(din_34_msk_ab0), .msk_a2b1(din_34_msk_ab1),
           .msk_a2b0_1sc(din_34_msk_ab0_1sc), .msk_a2b1_1sc(din_34_msk_ab1_1sc),
           
           .a3b0(din_36_ab0),
           .a3b0_1sc(din_36_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12)
) addr_5_31_calc (
           .clk(clk), .sign(din_signs_reg[31]), 
           .p(addr_5_31),
           .a0b0(din_31_ab0), .a0b1(din_31_ab1), .a0b2(din_31_ab2), .a0b3(din_31_ab3),
           .a0b0_1sc(din_31_ab0_1sc), .a0b1_1sc(din_31_ab1_1sc), .a0b2_1sc(din_31_ab2_1sc), .a0b3_1sc(din_31_ab3_1sc),
           .msk_a0b0(din_31_msk_ab0), .msk_a0b1(din_31_msk_ab1), .msk_a0b2(din_31_msk_ab2), .msk_a0b3(din_31_msk_ab3),
           .msk_a0b0_1sc(din_31_msk_ab0_1sc), .msk_a0b1_1sc(din_31_msk_ab1_1sc), .msk_a0b2_1sc(din_31_msk_ab2_1sc), .msk_a0b3_1sc(din_31_msk_ab3_1sc),

           .a1b0(din_33_ab0), .a1b1(din_33_ab1), .a1b2(din_33_ab2),
           .a1b0_1sc(din_33_ab0_1sc), .a1b1_1sc(din_33_ab1_1sc), .a1b2_1sc(din_33_ab2_1sc),
           .msk_a1b0(din_33_msk_ab0), .msk_a1b1(din_33_msk_ab1), .msk_a1b2(din_33_msk_ab2),
           .msk_a1b0_1sc(din_33_msk_ab0_1sc), .msk_a1b1_1sc(din_33_msk_ab1_1sc), .msk_a1b2_1sc(din_33_msk_ab2_1sc),

           .a2b0(din_35_ab0), .a2b1(din_35_ab1),
           .a2b0_1sc(din_35_ab0_1sc), .a2b1_1sc(din_35_ab1_1sc),
           .msk_a2b0(din_35_msk_ab0), .msk_a2b1(din_35_msk_ab1),
           .msk_a2b0_1sc(din_35_msk_ab0_1sc), .msk_a2b1_1sc(din_35_msk_ab1_1sc),
           
           .a3b0(din_37_ab0),
           .a3b0_1sc(din_37_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_0_calc (
           .clk(clk), .sign(din_signs_reg[0]), 
           .p(addr_6_0),
           .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
           .a0b0_1sc(din_0_ab0_1sc), .a0b1_1sc(din_0_ab1_1sc), .a0b2_1sc(din_0_ab2_1sc), .a0b3_1sc(din_0_ab3_1sc),
           .msk_a0b0(din_0_msk_ab0), .msk_a0b1(din_0_msk_ab1), .msk_a0b2(din_0_msk_ab2), .msk_a0b3(din_0_msk_ab3),
           .msk_a0b0_1sc(din_0_msk_ab0_1sc), .msk_a0b1_1sc(din_0_msk_ab1_1sc), .msk_a0b2_1sc(din_0_msk_ab2_1sc), .msk_a0b3_1sc(din_0_msk_ab3_1sc),

           .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2),
           .a1b0_1sc(din_2_ab0_1sc), .a1b1_1sc(din_2_ab1_1sc), .a1b2_1sc(din_2_ab2_1sc),
           .msk_a1b0(din_2_msk_ab0), .msk_a1b1(din_2_msk_ab1), .msk_a1b2(din_2_msk_ab2),
           .msk_a1b0_1sc(din_2_msk_ab0_1sc), .msk_a1b1_1sc(din_2_msk_ab1_1sc), .msk_a1b2_1sc(din_2_msk_ab2_1sc),

           .a2b0(din_4_ab0), .a2b1(din_4_ab1),
           .a2b0_1sc(din_4_ab0_1sc), .a2b1_1sc(din_4_ab1_1sc),
           .msk_a2b0(din_4_msk_ab0), .msk_a2b1(din_4_msk_ab1),
           .msk_a2b0_1sc(din_4_msk_ab0_1sc), .msk_a2b1_1sc(din_4_msk_ab1_1sc),
           
           .a3b0(din_6_ab0),
           .a3b0_1sc(din_6_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_1_calc (
           .clk(clk), .sign(din_signs_reg[1]), 
           .p(addr_6_1),
           .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
           .a0b0_1sc(din_1_ab0_1sc), .a0b1_1sc(din_1_ab1_1sc), .a0b2_1sc(din_1_ab2_1sc), .a0b3_1sc(din_1_ab3_1sc),
           .msk_a0b0(din_1_msk_ab0), .msk_a0b1(din_1_msk_ab1), .msk_a0b2(din_1_msk_ab2), .msk_a0b3(din_1_msk_ab3),
           .msk_a0b0_1sc(din_1_msk_ab0_1sc), .msk_a0b1_1sc(din_1_msk_ab1_1sc), .msk_a0b2_1sc(din_1_msk_ab2_1sc), .msk_a0b3_1sc(din_1_msk_ab3_1sc),

           .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2),
           .a1b0_1sc(din_3_ab0_1sc), .a1b1_1sc(din_3_ab1_1sc), .a1b2_1sc(din_3_ab2_1sc),
           .msk_a1b0(din_3_msk_ab0), .msk_a1b1(din_3_msk_ab1), .msk_a1b2(din_3_msk_ab2),
           .msk_a1b0_1sc(din_3_msk_ab0_1sc), .msk_a1b1_1sc(din_3_msk_ab1_1sc), .msk_a1b2_1sc(din_3_msk_ab2_1sc),

           .a2b0(din_5_ab0), .a2b1(din_5_ab1),
           .a2b0_1sc(din_5_ab0_1sc), .a2b1_1sc(din_5_ab1_1sc),
           .msk_a2b0(din_5_msk_ab0), .msk_a2b1(din_5_msk_ab1),
           .msk_a2b0_1sc(din_5_msk_ab0_1sc), .msk_a2b1_1sc(din_5_msk_ab1_1sc),
           
           .a3b0(din_7_ab0),
           .a3b0_1sc(din_7_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_2_calc (
           .clk(clk), .sign(din_signs_reg[2]), 
           .p(addr_6_2),
           .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
           .a0b0_1sc(din_2_ab0_1sc), .a0b1_1sc(din_2_ab1_1sc), .a0b2_1sc(din_2_ab2_1sc), .a0b3_1sc(din_2_ab3_1sc),
           .msk_a0b0(din_2_msk_ab0), .msk_a0b1(din_2_msk_ab1), .msk_a0b2(din_2_msk_ab2), .msk_a0b3(din_2_msk_ab3),
           .msk_a0b0_1sc(din_2_msk_ab0_1sc), .msk_a0b1_1sc(din_2_msk_ab1_1sc), .msk_a0b2_1sc(din_2_msk_ab2_1sc), .msk_a0b3_1sc(din_2_msk_ab3_1sc),

           .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2),
           .a1b0_1sc(din_4_ab0_1sc), .a1b1_1sc(din_4_ab1_1sc), .a1b2_1sc(din_4_ab2_1sc),
           .msk_a1b0(din_4_msk_ab0), .msk_a1b1(din_4_msk_ab1), .msk_a1b2(din_4_msk_ab2),
           .msk_a1b0_1sc(din_4_msk_ab0_1sc), .msk_a1b1_1sc(din_4_msk_ab1_1sc), .msk_a1b2_1sc(din_4_msk_ab2_1sc),

           .a2b0(din_6_ab0), .a2b1(din_6_ab1),
           .a2b0_1sc(din_6_ab0_1sc), .a2b1_1sc(din_6_ab1_1sc),
           .msk_a2b0(din_6_msk_ab0), .msk_a2b1(din_6_msk_ab1),
           .msk_a2b0_1sc(din_6_msk_ab0_1sc), .msk_a2b1_1sc(din_6_msk_ab1_1sc),
           
           .a3b0(din_8_ab0),
           .a3b0_1sc(din_8_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_3_calc (
           .clk(clk), .sign(din_signs_reg[3]), 
           .p(addr_6_3),
           .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
           .a0b0_1sc(din_3_ab0_1sc), .a0b1_1sc(din_3_ab1_1sc), .a0b2_1sc(din_3_ab2_1sc), .a0b3_1sc(din_3_ab3_1sc),
           .msk_a0b0(din_3_msk_ab0), .msk_a0b1(din_3_msk_ab1), .msk_a0b2(din_3_msk_ab2), .msk_a0b3(din_3_msk_ab3),
           .msk_a0b0_1sc(din_3_msk_ab0_1sc), .msk_a0b1_1sc(din_3_msk_ab1_1sc), .msk_a0b2_1sc(din_3_msk_ab2_1sc), .msk_a0b3_1sc(din_3_msk_ab3_1sc),

           .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2),
           .a1b0_1sc(din_5_ab0_1sc), .a1b1_1sc(din_5_ab1_1sc), .a1b2_1sc(din_5_ab2_1sc),
           .msk_a1b0(din_5_msk_ab0), .msk_a1b1(din_5_msk_ab1), .msk_a1b2(din_5_msk_ab2),
           .msk_a1b0_1sc(din_5_msk_ab0_1sc), .msk_a1b1_1sc(din_5_msk_ab1_1sc), .msk_a1b2_1sc(din_5_msk_ab2_1sc),

           .a2b0(din_7_ab0), .a2b1(din_7_ab1),
           .a2b0_1sc(din_7_ab0_1sc), .a2b1_1sc(din_7_ab1_1sc),
           .msk_a2b0(din_7_msk_ab0), .msk_a2b1(din_7_msk_ab1),
           .msk_a2b0_1sc(din_7_msk_ab0_1sc), .msk_a2b1_1sc(din_7_msk_ab1_1sc),
           
           .a3b0(din_9_ab0),
           .a3b0_1sc(din_9_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_4_calc (
           .clk(clk), .sign(din_signs_reg[4]), 
           .p(addr_6_4),
           .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
           .a0b0_1sc(din_4_ab0_1sc), .a0b1_1sc(din_4_ab1_1sc), .a0b2_1sc(din_4_ab2_1sc), .a0b3_1sc(din_4_ab3_1sc),
           .msk_a0b0(din_4_msk_ab0), .msk_a0b1(din_4_msk_ab1), .msk_a0b2(din_4_msk_ab2), .msk_a0b3(din_4_msk_ab3),
           .msk_a0b0_1sc(din_4_msk_ab0_1sc), .msk_a0b1_1sc(din_4_msk_ab1_1sc), .msk_a0b2_1sc(din_4_msk_ab2_1sc), .msk_a0b3_1sc(din_4_msk_ab3_1sc),

           .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2),
           .a1b0_1sc(din_6_ab0_1sc), .a1b1_1sc(din_6_ab1_1sc), .a1b2_1sc(din_6_ab2_1sc),
           .msk_a1b0(din_6_msk_ab0), .msk_a1b1(din_6_msk_ab1), .msk_a1b2(din_6_msk_ab2),
           .msk_a1b0_1sc(din_6_msk_ab0_1sc), .msk_a1b1_1sc(din_6_msk_ab1_1sc), .msk_a1b2_1sc(din_6_msk_ab2_1sc),

           .a2b0(din_8_ab0), .a2b1(din_8_ab1),
           .a2b0_1sc(din_8_ab0_1sc), .a2b1_1sc(din_8_ab1_1sc),
           .msk_a2b0(din_8_msk_ab0), .msk_a2b1(din_8_msk_ab1),
           .msk_a2b0_1sc(din_8_msk_ab0_1sc), .msk_a2b1_1sc(din_8_msk_ab1_1sc),
           
           .a3b0(din_10_ab0),
           .a3b0_1sc(din_10_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_5_calc (
           .clk(clk), .sign(din_signs_reg[5]), 
           .p(addr_6_5),
           .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
           .a0b0_1sc(din_5_ab0_1sc), .a0b1_1sc(din_5_ab1_1sc), .a0b2_1sc(din_5_ab2_1sc), .a0b3_1sc(din_5_ab3_1sc),
           .msk_a0b0(din_5_msk_ab0), .msk_a0b1(din_5_msk_ab1), .msk_a0b2(din_5_msk_ab2), .msk_a0b3(din_5_msk_ab3),
           .msk_a0b0_1sc(din_5_msk_ab0_1sc), .msk_a0b1_1sc(din_5_msk_ab1_1sc), .msk_a0b2_1sc(din_5_msk_ab2_1sc), .msk_a0b3_1sc(din_5_msk_ab3_1sc),

           .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2),
           .a1b0_1sc(din_7_ab0_1sc), .a1b1_1sc(din_7_ab1_1sc), .a1b2_1sc(din_7_ab2_1sc),
           .msk_a1b0(din_7_msk_ab0), .msk_a1b1(din_7_msk_ab1), .msk_a1b2(din_7_msk_ab2),
           .msk_a1b0_1sc(din_7_msk_ab0_1sc), .msk_a1b1_1sc(din_7_msk_ab1_1sc), .msk_a1b2_1sc(din_7_msk_ab2_1sc),

           .a2b0(din_9_ab0), .a2b1(din_9_ab1),
           .a2b0_1sc(din_9_ab0_1sc), .a2b1_1sc(din_9_ab1_1sc),
           .msk_a2b0(din_9_msk_ab0), .msk_a2b1(din_9_msk_ab1),
           .msk_a2b0_1sc(din_9_msk_ab0_1sc), .msk_a2b1_1sc(din_9_msk_ab1_1sc),
           
           .a3b0(din_11_ab0),
           .a3b0_1sc(din_11_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_6_calc (
           .clk(clk), .sign(din_signs_reg[6]), 
           .p(addr_6_6),
           .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
           .a0b0_1sc(din_6_ab0_1sc), .a0b1_1sc(din_6_ab1_1sc), .a0b2_1sc(din_6_ab2_1sc), .a0b3_1sc(din_6_ab3_1sc),
           .msk_a0b0(din_6_msk_ab0), .msk_a0b1(din_6_msk_ab1), .msk_a0b2(din_6_msk_ab2), .msk_a0b3(din_6_msk_ab3),
           .msk_a0b0_1sc(din_6_msk_ab0_1sc), .msk_a0b1_1sc(din_6_msk_ab1_1sc), .msk_a0b2_1sc(din_6_msk_ab2_1sc), .msk_a0b3_1sc(din_6_msk_ab3_1sc),

           .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2),
           .a1b0_1sc(din_8_ab0_1sc), .a1b1_1sc(din_8_ab1_1sc), .a1b2_1sc(din_8_ab2_1sc),
           .msk_a1b0(din_8_msk_ab0), .msk_a1b1(din_8_msk_ab1), .msk_a1b2(din_8_msk_ab2),
           .msk_a1b0_1sc(din_8_msk_ab0_1sc), .msk_a1b1_1sc(din_8_msk_ab1_1sc), .msk_a1b2_1sc(din_8_msk_ab2_1sc),

           .a2b0(din_10_ab0), .a2b1(din_10_ab1),
           .a2b0_1sc(din_10_ab0_1sc), .a2b1_1sc(din_10_ab1_1sc),
           .msk_a2b0(din_10_msk_ab0), .msk_a2b1(din_10_msk_ab1),
           .msk_a2b0_1sc(din_10_msk_ab0_1sc), .msk_a2b1_1sc(din_10_msk_ab1_1sc),
           
           .a3b0(din_12_ab0),
           .a3b0_1sc(din_12_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_7_calc (
           .clk(clk), .sign(din_signs_reg[7]), 
           .p(addr_6_7),
           .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
           .a0b0_1sc(din_7_ab0_1sc), .a0b1_1sc(din_7_ab1_1sc), .a0b2_1sc(din_7_ab2_1sc), .a0b3_1sc(din_7_ab3_1sc),
           .msk_a0b0(din_7_msk_ab0), .msk_a0b1(din_7_msk_ab1), .msk_a0b2(din_7_msk_ab2), .msk_a0b3(din_7_msk_ab3),
           .msk_a0b0_1sc(din_7_msk_ab0_1sc), .msk_a0b1_1sc(din_7_msk_ab1_1sc), .msk_a0b2_1sc(din_7_msk_ab2_1sc), .msk_a0b3_1sc(din_7_msk_ab3_1sc),

           .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2),
           .a1b0_1sc(din_9_ab0_1sc), .a1b1_1sc(din_9_ab1_1sc), .a1b2_1sc(din_9_ab2_1sc),
           .msk_a1b0(din_9_msk_ab0), .msk_a1b1(din_9_msk_ab1), .msk_a1b2(din_9_msk_ab2),
           .msk_a1b0_1sc(din_9_msk_ab0_1sc), .msk_a1b1_1sc(din_9_msk_ab1_1sc), .msk_a1b2_1sc(din_9_msk_ab2_1sc),

           .a2b0(din_11_ab0), .a2b1(din_11_ab1),
           .a2b0_1sc(din_11_ab0_1sc), .a2b1_1sc(din_11_ab1_1sc),
           .msk_a2b0(din_11_msk_ab0), .msk_a2b1(din_11_msk_ab1),
           .msk_a2b0_1sc(din_11_msk_ab0_1sc), .msk_a2b1_1sc(din_11_msk_ab1_1sc),
           
           .a3b0(din_13_ab0),
           .a3b0_1sc(din_13_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_8_calc (
           .clk(clk), .sign(din_signs_reg[8]), 
           .p(addr_6_8),
           .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
           .a0b0_1sc(din_8_ab0_1sc), .a0b1_1sc(din_8_ab1_1sc), .a0b2_1sc(din_8_ab2_1sc), .a0b3_1sc(din_8_ab3_1sc),
           .msk_a0b0(din_8_msk_ab0), .msk_a0b1(din_8_msk_ab1), .msk_a0b2(din_8_msk_ab2), .msk_a0b3(din_8_msk_ab3),
           .msk_a0b0_1sc(din_8_msk_ab0_1sc), .msk_a0b1_1sc(din_8_msk_ab1_1sc), .msk_a0b2_1sc(din_8_msk_ab2_1sc), .msk_a0b3_1sc(din_8_msk_ab3_1sc),

           .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2),
           .a1b0_1sc(din_10_ab0_1sc), .a1b1_1sc(din_10_ab1_1sc), .a1b2_1sc(din_10_ab2_1sc),
           .msk_a1b0(din_10_msk_ab0), .msk_a1b1(din_10_msk_ab1), .msk_a1b2(din_10_msk_ab2),
           .msk_a1b0_1sc(din_10_msk_ab0_1sc), .msk_a1b1_1sc(din_10_msk_ab1_1sc), .msk_a1b2_1sc(din_10_msk_ab2_1sc),

           .a2b0(din_12_ab0), .a2b1(din_12_ab1),
           .a2b0_1sc(din_12_ab0_1sc), .a2b1_1sc(din_12_ab1_1sc),
           .msk_a2b0(din_12_msk_ab0), .msk_a2b1(din_12_msk_ab1),
           .msk_a2b0_1sc(din_12_msk_ab0_1sc), .msk_a2b1_1sc(din_12_msk_ab1_1sc),
           
           .a3b0(din_14_ab0),
           .a3b0_1sc(din_14_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_9_calc (
           .clk(clk), .sign(din_signs_reg[9]), 
           .p(addr_6_9),
           .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
           .a0b0_1sc(din_9_ab0_1sc), .a0b1_1sc(din_9_ab1_1sc), .a0b2_1sc(din_9_ab2_1sc), .a0b3_1sc(din_9_ab3_1sc),
           .msk_a0b0(din_9_msk_ab0), .msk_a0b1(din_9_msk_ab1), .msk_a0b2(din_9_msk_ab2), .msk_a0b3(din_9_msk_ab3),
           .msk_a0b0_1sc(din_9_msk_ab0_1sc), .msk_a0b1_1sc(din_9_msk_ab1_1sc), .msk_a0b2_1sc(din_9_msk_ab2_1sc), .msk_a0b3_1sc(din_9_msk_ab3_1sc),

           .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2),
           .a1b0_1sc(din_11_ab0_1sc), .a1b1_1sc(din_11_ab1_1sc), .a1b2_1sc(din_11_ab2_1sc),
           .msk_a1b0(din_11_msk_ab0), .msk_a1b1(din_11_msk_ab1), .msk_a1b2(din_11_msk_ab2),
           .msk_a1b0_1sc(din_11_msk_ab0_1sc), .msk_a1b1_1sc(din_11_msk_ab1_1sc), .msk_a1b2_1sc(din_11_msk_ab2_1sc),

           .a2b0(din_13_ab0), .a2b1(din_13_ab1),
           .a2b0_1sc(din_13_ab0_1sc), .a2b1_1sc(din_13_ab1_1sc),
           .msk_a2b0(din_13_msk_ab0), .msk_a2b1(din_13_msk_ab1),
           .msk_a2b0_1sc(din_13_msk_ab0_1sc), .msk_a2b1_1sc(din_13_msk_ab1_1sc),
           
           .a3b0(din_15_ab0),
           .a3b0_1sc(din_15_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_10_calc (
           .clk(clk), .sign(din_signs_reg[10]), 
           .p(addr_6_10),
           .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
           .a0b0_1sc(din_10_ab0_1sc), .a0b1_1sc(din_10_ab1_1sc), .a0b2_1sc(din_10_ab2_1sc), .a0b3_1sc(din_10_ab3_1sc),
           .msk_a0b0(din_10_msk_ab0), .msk_a0b1(din_10_msk_ab1), .msk_a0b2(din_10_msk_ab2), .msk_a0b3(din_10_msk_ab3),
           .msk_a0b0_1sc(din_10_msk_ab0_1sc), .msk_a0b1_1sc(din_10_msk_ab1_1sc), .msk_a0b2_1sc(din_10_msk_ab2_1sc), .msk_a0b3_1sc(din_10_msk_ab3_1sc),

           .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2),
           .a1b0_1sc(din_12_ab0_1sc), .a1b1_1sc(din_12_ab1_1sc), .a1b2_1sc(din_12_ab2_1sc),
           .msk_a1b0(din_12_msk_ab0), .msk_a1b1(din_12_msk_ab1), .msk_a1b2(din_12_msk_ab2),
           .msk_a1b0_1sc(din_12_msk_ab0_1sc), .msk_a1b1_1sc(din_12_msk_ab1_1sc), .msk_a1b2_1sc(din_12_msk_ab2_1sc),

           .a2b0(din_14_ab0), .a2b1(din_14_ab1),
           .a2b0_1sc(din_14_ab0_1sc), .a2b1_1sc(din_14_ab1_1sc),
           .msk_a2b0(din_14_msk_ab0), .msk_a2b1(din_14_msk_ab1),
           .msk_a2b0_1sc(din_14_msk_ab0_1sc), .msk_a2b1_1sc(din_14_msk_ab1_1sc),
           
           .a3b0(din_16_ab0),
           .a3b0_1sc(din_16_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_11_calc (
           .clk(clk), .sign(din_signs_reg[11]), 
           .p(addr_6_11),
           .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
           .a0b0_1sc(din_11_ab0_1sc), .a0b1_1sc(din_11_ab1_1sc), .a0b2_1sc(din_11_ab2_1sc), .a0b3_1sc(din_11_ab3_1sc),
           .msk_a0b0(din_11_msk_ab0), .msk_a0b1(din_11_msk_ab1), .msk_a0b2(din_11_msk_ab2), .msk_a0b3(din_11_msk_ab3),
           .msk_a0b0_1sc(din_11_msk_ab0_1sc), .msk_a0b1_1sc(din_11_msk_ab1_1sc), .msk_a0b2_1sc(din_11_msk_ab2_1sc), .msk_a0b3_1sc(din_11_msk_ab3_1sc),

           .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2),
           .a1b0_1sc(din_13_ab0_1sc), .a1b1_1sc(din_13_ab1_1sc), .a1b2_1sc(din_13_ab2_1sc),
           .msk_a1b0(din_13_msk_ab0), .msk_a1b1(din_13_msk_ab1), .msk_a1b2(din_13_msk_ab2),
           .msk_a1b0_1sc(din_13_msk_ab0_1sc), .msk_a1b1_1sc(din_13_msk_ab1_1sc), .msk_a1b2_1sc(din_13_msk_ab2_1sc),

           .a2b0(din_15_ab0), .a2b1(din_15_ab1),
           .a2b0_1sc(din_15_ab0_1sc), .a2b1_1sc(din_15_ab1_1sc),
           .msk_a2b0(din_15_msk_ab0), .msk_a2b1(din_15_msk_ab1),
           .msk_a2b0_1sc(din_15_msk_ab0_1sc), .msk_a2b1_1sc(din_15_msk_ab1_1sc),
           
           .a3b0(din_17_ab0),
           .a3b0_1sc(din_17_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_12_calc (
           .clk(clk), .sign(din_signs_reg[12]), 
           .p(addr_6_12),
           .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
           .a0b0_1sc(din_12_ab0_1sc), .a0b1_1sc(din_12_ab1_1sc), .a0b2_1sc(din_12_ab2_1sc), .a0b3_1sc(din_12_ab3_1sc),
           .msk_a0b0(din_12_msk_ab0), .msk_a0b1(din_12_msk_ab1), .msk_a0b2(din_12_msk_ab2), .msk_a0b3(din_12_msk_ab3),
           .msk_a0b0_1sc(din_12_msk_ab0_1sc), .msk_a0b1_1sc(din_12_msk_ab1_1sc), .msk_a0b2_1sc(din_12_msk_ab2_1sc), .msk_a0b3_1sc(din_12_msk_ab3_1sc),

           .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2),
           .a1b0_1sc(din_14_ab0_1sc), .a1b1_1sc(din_14_ab1_1sc), .a1b2_1sc(din_14_ab2_1sc),
           .msk_a1b0(din_14_msk_ab0), .msk_a1b1(din_14_msk_ab1), .msk_a1b2(din_14_msk_ab2),
           .msk_a1b0_1sc(din_14_msk_ab0_1sc), .msk_a1b1_1sc(din_14_msk_ab1_1sc), .msk_a1b2_1sc(din_14_msk_ab2_1sc),

           .a2b0(din_16_ab0), .a2b1(din_16_ab1),
           .a2b0_1sc(din_16_ab0_1sc), .a2b1_1sc(din_16_ab1_1sc),
           .msk_a2b0(din_16_msk_ab0), .msk_a2b1(din_16_msk_ab1),
           .msk_a2b0_1sc(din_16_msk_ab0_1sc), .msk_a2b1_1sc(din_16_msk_ab1_1sc),
           
           .a3b0(din_18_ab0),
           .a3b0_1sc(din_18_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_13_calc (
           .clk(clk), .sign(din_signs_reg[13]), 
           .p(addr_6_13),
           .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
           .a0b0_1sc(din_13_ab0_1sc), .a0b1_1sc(din_13_ab1_1sc), .a0b2_1sc(din_13_ab2_1sc), .a0b3_1sc(din_13_ab3_1sc),
           .msk_a0b0(din_13_msk_ab0), .msk_a0b1(din_13_msk_ab1), .msk_a0b2(din_13_msk_ab2), .msk_a0b3(din_13_msk_ab3),
           .msk_a0b0_1sc(din_13_msk_ab0_1sc), .msk_a0b1_1sc(din_13_msk_ab1_1sc), .msk_a0b2_1sc(din_13_msk_ab2_1sc), .msk_a0b3_1sc(din_13_msk_ab3_1sc),

           .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2),
           .a1b0_1sc(din_15_ab0_1sc), .a1b1_1sc(din_15_ab1_1sc), .a1b2_1sc(din_15_ab2_1sc),
           .msk_a1b0(din_15_msk_ab0), .msk_a1b1(din_15_msk_ab1), .msk_a1b2(din_15_msk_ab2),
           .msk_a1b0_1sc(din_15_msk_ab0_1sc), .msk_a1b1_1sc(din_15_msk_ab1_1sc), .msk_a1b2_1sc(din_15_msk_ab2_1sc),

           .a2b0(din_17_ab0), .a2b1(din_17_ab1),
           .a2b0_1sc(din_17_ab0_1sc), .a2b1_1sc(din_17_ab1_1sc),
           .msk_a2b0(din_17_msk_ab0), .msk_a2b1(din_17_msk_ab1),
           .msk_a2b0_1sc(din_17_msk_ab0_1sc), .msk_a2b1_1sc(din_17_msk_ab1_1sc),
           
           .a3b0(din_19_ab0),
           .a3b0_1sc(din_19_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_14_calc (
           .clk(clk), .sign(din_signs_reg[14]), 
           .p(addr_6_14),
           .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
           .a0b0_1sc(din_14_ab0_1sc), .a0b1_1sc(din_14_ab1_1sc), .a0b2_1sc(din_14_ab2_1sc), .a0b3_1sc(din_14_ab3_1sc),
           .msk_a0b0(din_14_msk_ab0), .msk_a0b1(din_14_msk_ab1), .msk_a0b2(din_14_msk_ab2), .msk_a0b3(din_14_msk_ab3),
           .msk_a0b0_1sc(din_14_msk_ab0_1sc), .msk_a0b1_1sc(din_14_msk_ab1_1sc), .msk_a0b2_1sc(din_14_msk_ab2_1sc), .msk_a0b3_1sc(din_14_msk_ab3_1sc),

           .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2),
           .a1b0_1sc(din_16_ab0_1sc), .a1b1_1sc(din_16_ab1_1sc), .a1b2_1sc(din_16_ab2_1sc),
           .msk_a1b0(din_16_msk_ab0), .msk_a1b1(din_16_msk_ab1), .msk_a1b2(din_16_msk_ab2),
           .msk_a1b0_1sc(din_16_msk_ab0_1sc), .msk_a1b1_1sc(din_16_msk_ab1_1sc), .msk_a1b2_1sc(din_16_msk_ab2_1sc),

           .a2b0(din_18_ab0), .a2b1(din_18_ab1),
           .a2b0_1sc(din_18_ab0_1sc), .a2b1_1sc(din_18_ab1_1sc),
           .msk_a2b0(din_18_msk_ab0), .msk_a2b1(din_18_msk_ab1),
           .msk_a2b0_1sc(din_18_msk_ab0_1sc), .msk_a2b1_1sc(din_18_msk_ab1_1sc),
           
           .a3b0(din_20_ab0),
           .a3b0_1sc(din_20_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_15_calc (
           .clk(clk), .sign(din_signs_reg[15]), 
           .p(addr_6_15),
           .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
           .a0b0_1sc(din_15_ab0_1sc), .a0b1_1sc(din_15_ab1_1sc), .a0b2_1sc(din_15_ab2_1sc), .a0b3_1sc(din_15_ab3_1sc),
           .msk_a0b0(din_15_msk_ab0), .msk_a0b1(din_15_msk_ab1), .msk_a0b2(din_15_msk_ab2), .msk_a0b3(din_15_msk_ab3),
           .msk_a0b0_1sc(din_15_msk_ab0_1sc), .msk_a0b1_1sc(din_15_msk_ab1_1sc), .msk_a0b2_1sc(din_15_msk_ab2_1sc), .msk_a0b3_1sc(din_15_msk_ab3_1sc),

           .a1b0(din_17_ab0), .a1b1(din_17_ab1), .a1b2(din_17_ab2),
           .a1b0_1sc(din_17_ab0_1sc), .a1b1_1sc(din_17_ab1_1sc), .a1b2_1sc(din_17_ab2_1sc),
           .msk_a1b0(din_17_msk_ab0), .msk_a1b1(din_17_msk_ab1), .msk_a1b2(din_17_msk_ab2),
           .msk_a1b0_1sc(din_17_msk_ab0_1sc), .msk_a1b1_1sc(din_17_msk_ab1_1sc), .msk_a1b2_1sc(din_17_msk_ab2_1sc),

           .a2b0(din_19_ab0), .a2b1(din_19_ab1),
           .a2b0_1sc(din_19_ab0_1sc), .a2b1_1sc(din_19_ab1_1sc),
           .msk_a2b0(din_19_msk_ab0), .msk_a2b1(din_19_msk_ab1),
           .msk_a2b0_1sc(din_19_msk_ab0_1sc), .msk_a2b1_1sc(din_19_msk_ab1_1sc),
           
           .a3b0(din_21_ab0),
           .a3b0_1sc(din_21_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_16_calc (
           .clk(clk), .sign(din_signs_reg[16]), 
           .p(addr_6_16),
           .a0b0(din_16_ab0), .a0b1(din_16_ab1), .a0b2(din_16_ab2), .a0b3(din_16_ab3),
           .a0b0_1sc(din_16_ab0_1sc), .a0b1_1sc(din_16_ab1_1sc), .a0b2_1sc(din_16_ab2_1sc), .a0b3_1sc(din_16_ab3_1sc),
           .msk_a0b0(din_16_msk_ab0), .msk_a0b1(din_16_msk_ab1), .msk_a0b2(din_16_msk_ab2), .msk_a0b3(din_16_msk_ab3),
           .msk_a0b0_1sc(din_16_msk_ab0_1sc), .msk_a0b1_1sc(din_16_msk_ab1_1sc), .msk_a0b2_1sc(din_16_msk_ab2_1sc), .msk_a0b3_1sc(din_16_msk_ab3_1sc),

           .a1b0(din_18_ab0), .a1b1(din_18_ab1), .a1b2(din_18_ab2),
           .a1b0_1sc(din_18_ab0_1sc), .a1b1_1sc(din_18_ab1_1sc), .a1b2_1sc(din_18_ab2_1sc),
           .msk_a1b0(din_18_msk_ab0), .msk_a1b1(din_18_msk_ab1), .msk_a1b2(din_18_msk_ab2),
           .msk_a1b0_1sc(din_18_msk_ab0_1sc), .msk_a1b1_1sc(din_18_msk_ab1_1sc), .msk_a1b2_1sc(din_18_msk_ab2_1sc),

           .a2b0(din_20_ab0), .a2b1(din_20_ab1),
           .a2b0_1sc(din_20_ab0_1sc), .a2b1_1sc(din_20_ab1_1sc),
           .msk_a2b0(din_20_msk_ab0), .msk_a2b1(din_20_msk_ab1),
           .msk_a2b0_1sc(din_20_msk_ab0_1sc), .msk_a2b1_1sc(din_20_msk_ab1_1sc),
           
           .a3b0(din_22_ab0),
           .a3b0_1sc(din_22_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_17_calc (
           .clk(clk), .sign(din_signs_reg[17]), 
           .p(addr_6_17),
           .a0b0(din_17_ab0), .a0b1(din_17_ab1), .a0b2(din_17_ab2), .a0b3(din_17_ab3),
           .a0b0_1sc(din_17_ab0_1sc), .a0b1_1sc(din_17_ab1_1sc), .a0b2_1sc(din_17_ab2_1sc), .a0b3_1sc(din_17_ab3_1sc),
           .msk_a0b0(din_17_msk_ab0), .msk_a0b1(din_17_msk_ab1), .msk_a0b2(din_17_msk_ab2), .msk_a0b3(din_17_msk_ab3),
           .msk_a0b0_1sc(din_17_msk_ab0_1sc), .msk_a0b1_1sc(din_17_msk_ab1_1sc), .msk_a0b2_1sc(din_17_msk_ab2_1sc), .msk_a0b3_1sc(din_17_msk_ab3_1sc),

           .a1b0(din_19_ab0), .a1b1(din_19_ab1), .a1b2(din_19_ab2),
           .a1b0_1sc(din_19_ab0_1sc), .a1b1_1sc(din_19_ab1_1sc), .a1b2_1sc(din_19_ab2_1sc),
           .msk_a1b0(din_19_msk_ab0), .msk_a1b1(din_19_msk_ab1), .msk_a1b2(din_19_msk_ab2),
           .msk_a1b0_1sc(din_19_msk_ab0_1sc), .msk_a1b1_1sc(din_19_msk_ab1_1sc), .msk_a1b2_1sc(din_19_msk_ab2_1sc),

           .a2b0(din_21_ab0), .a2b1(din_21_ab1),
           .a2b0_1sc(din_21_ab0_1sc), .a2b1_1sc(din_21_ab1_1sc),
           .msk_a2b0(din_21_msk_ab0), .msk_a2b1(din_21_msk_ab1),
           .msk_a2b0_1sc(din_21_msk_ab0_1sc), .msk_a2b1_1sc(din_21_msk_ab1_1sc),
           
           .a3b0(din_23_ab0),
           .a3b0_1sc(din_23_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_18_calc (
           .clk(clk), .sign(din_signs_reg[18]), 
           .p(addr_6_18),
           .a0b0(din_18_ab0), .a0b1(din_18_ab1), .a0b2(din_18_ab2), .a0b3(din_18_ab3),
           .a0b0_1sc(din_18_ab0_1sc), .a0b1_1sc(din_18_ab1_1sc), .a0b2_1sc(din_18_ab2_1sc), .a0b3_1sc(din_18_ab3_1sc),
           .msk_a0b0(din_18_msk_ab0), .msk_a0b1(din_18_msk_ab1), .msk_a0b2(din_18_msk_ab2), .msk_a0b3(din_18_msk_ab3),
           .msk_a0b0_1sc(din_18_msk_ab0_1sc), .msk_a0b1_1sc(din_18_msk_ab1_1sc), .msk_a0b2_1sc(din_18_msk_ab2_1sc), .msk_a0b3_1sc(din_18_msk_ab3_1sc),

           .a1b0(din_20_ab0), .a1b1(din_20_ab1), .a1b2(din_20_ab2),
           .a1b0_1sc(din_20_ab0_1sc), .a1b1_1sc(din_20_ab1_1sc), .a1b2_1sc(din_20_ab2_1sc),
           .msk_a1b0(din_20_msk_ab0), .msk_a1b1(din_20_msk_ab1), .msk_a1b2(din_20_msk_ab2),
           .msk_a1b0_1sc(din_20_msk_ab0_1sc), .msk_a1b1_1sc(din_20_msk_ab1_1sc), .msk_a1b2_1sc(din_20_msk_ab2_1sc),

           .a2b0(din_22_ab0), .a2b1(din_22_ab1),
           .a2b0_1sc(din_22_ab0_1sc), .a2b1_1sc(din_22_ab1_1sc),
           .msk_a2b0(din_22_msk_ab0), .msk_a2b1(din_22_msk_ab1),
           .msk_a2b0_1sc(din_22_msk_ab0_1sc), .msk_a2b1_1sc(din_22_msk_ab1_1sc),
           
           .a3b0(din_24_ab0),
           .a3b0_1sc(din_24_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_19_calc (
           .clk(clk), .sign(din_signs_reg[19]), 
           .p(addr_6_19),
           .a0b0(din_19_ab0), .a0b1(din_19_ab1), .a0b2(din_19_ab2), .a0b3(din_19_ab3),
           .a0b0_1sc(din_19_ab0_1sc), .a0b1_1sc(din_19_ab1_1sc), .a0b2_1sc(din_19_ab2_1sc), .a0b3_1sc(din_19_ab3_1sc),
           .msk_a0b0(din_19_msk_ab0), .msk_a0b1(din_19_msk_ab1), .msk_a0b2(din_19_msk_ab2), .msk_a0b3(din_19_msk_ab3),
           .msk_a0b0_1sc(din_19_msk_ab0_1sc), .msk_a0b1_1sc(din_19_msk_ab1_1sc), .msk_a0b2_1sc(din_19_msk_ab2_1sc), .msk_a0b3_1sc(din_19_msk_ab3_1sc),

           .a1b0(din_21_ab0), .a1b1(din_21_ab1), .a1b2(din_21_ab2),
           .a1b0_1sc(din_21_ab0_1sc), .a1b1_1sc(din_21_ab1_1sc), .a1b2_1sc(din_21_ab2_1sc),
           .msk_a1b0(din_21_msk_ab0), .msk_a1b1(din_21_msk_ab1), .msk_a1b2(din_21_msk_ab2),
           .msk_a1b0_1sc(din_21_msk_ab0_1sc), .msk_a1b1_1sc(din_21_msk_ab1_1sc), .msk_a1b2_1sc(din_21_msk_ab2_1sc),

           .a2b0(din_23_ab0), .a2b1(din_23_ab1),
           .a2b0_1sc(din_23_ab0_1sc), .a2b1_1sc(din_23_ab1_1sc),
           .msk_a2b0(din_23_msk_ab0), .msk_a2b1(din_23_msk_ab1),
           .msk_a2b0_1sc(din_23_msk_ab0_1sc), .msk_a2b1_1sc(din_23_msk_ab1_1sc),
           
           .a3b0(din_25_ab0),
           .a3b0_1sc(din_25_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_20_calc (
           .clk(clk), .sign(din_signs_reg[20]), 
           .p(addr_6_20),
           .a0b0(din_20_ab0), .a0b1(din_20_ab1), .a0b2(din_20_ab2), .a0b3(din_20_ab3),
           .a0b0_1sc(din_20_ab0_1sc), .a0b1_1sc(din_20_ab1_1sc), .a0b2_1sc(din_20_ab2_1sc), .a0b3_1sc(din_20_ab3_1sc),
           .msk_a0b0(din_20_msk_ab0), .msk_a0b1(din_20_msk_ab1), .msk_a0b2(din_20_msk_ab2), .msk_a0b3(din_20_msk_ab3),
           .msk_a0b0_1sc(din_20_msk_ab0_1sc), .msk_a0b1_1sc(din_20_msk_ab1_1sc), .msk_a0b2_1sc(din_20_msk_ab2_1sc), .msk_a0b3_1sc(din_20_msk_ab3_1sc),

           .a1b0(din_22_ab0), .a1b1(din_22_ab1), .a1b2(din_22_ab2),
           .a1b0_1sc(din_22_ab0_1sc), .a1b1_1sc(din_22_ab1_1sc), .a1b2_1sc(din_22_ab2_1sc),
           .msk_a1b0(din_22_msk_ab0), .msk_a1b1(din_22_msk_ab1), .msk_a1b2(din_22_msk_ab2),
           .msk_a1b0_1sc(din_22_msk_ab0_1sc), .msk_a1b1_1sc(din_22_msk_ab1_1sc), .msk_a1b2_1sc(din_22_msk_ab2_1sc),

           .a2b0(din_24_ab0), .a2b1(din_24_ab1),
           .a2b0_1sc(din_24_ab0_1sc), .a2b1_1sc(din_24_ab1_1sc),
           .msk_a2b0(din_24_msk_ab0), .msk_a2b1(din_24_msk_ab1),
           .msk_a2b0_1sc(din_24_msk_ab0_1sc), .msk_a2b1_1sc(din_24_msk_ab1_1sc),
           
           .a3b0(din_26_ab0),
           .a3b0_1sc(din_26_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_21_calc (
           .clk(clk), .sign(din_signs_reg[21]), 
           .p(addr_6_21),
           .a0b0(din_21_ab0), .a0b1(din_21_ab1), .a0b2(din_21_ab2), .a0b3(din_21_ab3),
           .a0b0_1sc(din_21_ab0_1sc), .a0b1_1sc(din_21_ab1_1sc), .a0b2_1sc(din_21_ab2_1sc), .a0b3_1sc(din_21_ab3_1sc),
           .msk_a0b0(din_21_msk_ab0), .msk_a0b1(din_21_msk_ab1), .msk_a0b2(din_21_msk_ab2), .msk_a0b3(din_21_msk_ab3),
           .msk_a0b0_1sc(din_21_msk_ab0_1sc), .msk_a0b1_1sc(din_21_msk_ab1_1sc), .msk_a0b2_1sc(din_21_msk_ab2_1sc), .msk_a0b3_1sc(din_21_msk_ab3_1sc),

           .a1b0(din_23_ab0), .a1b1(din_23_ab1), .a1b2(din_23_ab2),
           .a1b0_1sc(din_23_ab0_1sc), .a1b1_1sc(din_23_ab1_1sc), .a1b2_1sc(din_23_ab2_1sc),
           .msk_a1b0(din_23_msk_ab0), .msk_a1b1(din_23_msk_ab1), .msk_a1b2(din_23_msk_ab2),
           .msk_a1b0_1sc(din_23_msk_ab0_1sc), .msk_a1b1_1sc(din_23_msk_ab1_1sc), .msk_a1b2_1sc(din_23_msk_ab2_1sc),

           .a2b0(din_25_ab0), .a2b1(din_25_ab1),
           .a2b0_1sc(din_25_ab0_1sc), .a2b1_1sc(din_25_ab1_1sc),
           .msk_a2b0(din_25_msk_ab0), .msk_a2b1(din_25_msk_ab1),
           .msk_a2b0_1sc(din_25_msk_ab0_1sc), .msk_a2b1_1sc(din_25_msk_ab1_1sc),
           
           .a3b0(din_27_ab0),
           .a3b0_1sc(din_27_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_22_calc (
           .clk(clk), .sign(din_signs_reg[22]), 
           .p(addr_6_22),
           .a0b0(din_22_ab0), .a0b1(din_22_ab1), .a0b2(din_22_ab2), .a0b3(din_22_ab3),
           .a0b0_1sc(din_22_ab0_1sc), .a0b1_1sc(din_22_ab1_1sc), .a0b2_1sc(din_22_ab2_1sc), .a0b3_1sc(din_22_ab3_1sc),
           .msk_a0b0(din_22_msk_ab0), .msk_a0b1(din_22_msk_ab1), .msk_a0b2(din_22_msk_ab2), .msk_a0b3(din_22_msk_ab3),
           .msk_a0b0_1sc(din_22_msk_ab0_1sc), .msk_a0b1_1sc(din_22_msk_ab1_1sc), .msk_a0b2_1sc(din_22_msk_ab2_1sc), .msk_a0b3_1sc(din_22_msk_ab3_1sc),

           .a1b0(din_24_ab0), .a1b1(din_24_ab1), .a1b2(din_24_ab2),
           .a1b0_1sc(din_24_ab0_1sc), .a1b1_1sc(din_24_ab1_1sc), .a1b2_1sc(din_24_ab2_1sc),
           .msk_a1b0(din_24_msk_ab0), .msk_a1b1(din_24_msk_ab1), .msk_a1b2(din_24_msk_ab2),
           .msk_a1b0_1sc(din_24_msk_ab0_1sc), .msk_a1b1_1sc(din_24_msk_ab1_1sc), .msk_a1b2_1sc(din_24_msk_ab2_1sc),

           .a2b0(din_26_ab0), .a2b1(din_26_ab1),
           .a2b0_1sc(din_26_ab0_1sc), .a2b1_1sc(din_26_ab1_1sc),
           .msk_a2b0(din_26_msk_ab0), .msk_a2b1(din_26_msk_ab1),
           .msk_a2b0_1sc(din_26_msk_ab0_1sc), .msk_a2b1_1sc(din_26_msk_ab1_1sc),
           
           .a3b0(din_28_ab0),
           .a3b0_1sc(din_28_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_23_calc (
           .clk(clk), .sign(din_signs_reg[23]), 
           .p(addr_6_23),
           .a0b0(din_23_ab0), .a0b1(din_23_ab1), .a0b2(din_23_ab2), .a0b3(din_23_ab3),
           .a0b0_1sc(din_23_ab0_1sc), .a0b1_1sc(din_23_ab1_1sc), .a0b2_1sc(din_23_ab2_1sc), .a0b3_1sc(din_23_ab3_1sc),
           .msk_a0b0(din_23_msk_ab0), .msk_a0b1(din_23_msk_ab1), .msk_a0b2(din_23_msk_ab2), .msk_a0b3(din_23_msk_ab3),
           .msk_a0b0_1sc(din_23_msk_ab0_1sc), .msk_a0b1_1sc(din_23_msk_ab1_1sc), .msk_a0b2_1sc(din_23_msk_ab2_1sc), .msk_a0b3_1sc(din_23_msk_ab3_1sc),

           .a1b0(din_25_ab0), .a1b1(din_25_ab1), .a1b2(din_25_ab2),
           .a1b0_1sc(din_25_ab0_1sc), .a1b1_1sc(din_25_ab1_1sc), .a1b2_1sc(din_25_ab2_1sc),
           .msk_a1b0(din_25_msk_ab0), .msk_a1b1(din_25_msk_ab1), .msk_a1b2(din_25_msk_ab2),
           .msk_a1b0_1sc(din_25_msk_ab0_1sc), .msk_a1b1_1sc(din_25_msk_ab1_1sc), .msk_a1b2_1sc(din_25_msk_ab2_1sc),

           .a2b0(din_27_ab0), .a2b1(din_27_ab1),
           .a2b0_1sc(din_27_ab0_1sc), .a2b1_1sc(din_27_ab1_1sc),
           .msk_a2b0(din_27_msk_ab0), .msk_a2b1(din_27_msk_ab1),
           .msk_a2b0_1sc(din_27_msk_ab0_1sc), .msk_a2b1_1sc(din_27_msk_ab1_1sc),
           
           .a3b0(din_29_ab0),
           .a3b0_1sc(din_29_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_24_calc (
           .clk(clk), .sign(din_signs_reg[24]), 
           .p(addr_6_24),
           .a0b0(din_24_ab0), .a0b1(din_24_ab1), .a0b2(din_24_ab2), .a0b3(din_24_ab3),
           .a0b0_1sc(din_24_ab0_1sc), .a0b1_1sc(din_24_ab1_1sc), .a0b2_1sc(din_24_ab2_1sc), .a0b3_1sc(din_24_ab3_1sc),
           .msk_a0b0(din_24_msk_ab0), .msk_a0b1(din_24_msk_ab1), .msk_a0b2(din_24_msk_ab2), .msk_a0b3(din_24_msk_ab3),
           .msk_a0b0_1sc(din_24_msk_ab0_1sc), .msk_a0b1_1sc(din_24_msk_ab1_1sc), .msk_a0b2_1sc(din_24_msk_ab2_1sc), .msk_a0b3_1sc(din_24_msk_ab3_1sc),

           .a1b0(din_26_ab0), .a1b1(din_26_ab1), .a1b2(din_26_ab2),
           .a1b0_1sc(din_26_ab0_1sc), .a1b1_1sc(din_26_ab1_1sc), .a1b2_1sc(din_26_ab2_1sc),
           .msk_a1b0(din_26_msk_ab0), .msk_a1b1(din_26_msk_ab1), .msk_a1b2(din_26_msk_ab2),
           .msk_a1b0_1sc(din_26_msk_ab0_1sc), .msk_a1b1_1sc(din_26_msk_ab1_1sc), .msk_a1b2_1sc(din_26_msk_ab2_1sc),

           .a2b0(din_28_ab0), .a2b1(din_28_ab1),
           .a2b0_1sc(din_28_ab0_1sc), .a2b1_1sc(din_28_ab1_1sc),
           .msk_a2b0(din_28_msk_ab0), .msk_a2b1(din_28_msk_ab1),
           .msk_a2b0_1sc(din_28_msk_ab0_1sc), .msk_a2b1_1sc(din_28_msk_ab1_1sc),
           
           .a3b0(din_30_ab0),
           .a3b0_1sc(din_30_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_25_calc (
           .clk(clk), .sign(din_signs_reg[25]), 
           .p(addr_6_25),
           .a0b0(din_25_ab0), .a0b1(din_25_ab1), .a0b2(din_25_ab2), .a0b3(din_25_ab3),
           .a0b0_1sc(din_25_ab0_1sc), .a0b1_1sc(din_25_ab1_1sc), .a0b2_1sc(din_25_ab2_1sc), .a0b3_1sc(din_25_ab3_1sc),
           .msk_a0b0(din_25_msk_ab0), .msk_a0b1(din_25_msk_ab1), .msk_a0b2(din_25_msk_ab2), .msk_a0b3(din_25_msk_ab3),
           .msk_a0b0_1sc(din_25_msk_ab0_1sc), .msk_a0b1_1sc(din_25_msk_ab1_1sc), .msk_a0b2_1sc(din_25_msk_ab2_1sc), .msk_a0b3_1sc(din_25_msk_ab3_1sc),

           .a1b0(din_27_ab0), .a1b1(din_27_ab1), .a1b2(din_27_ab2),
           .a1b0_1sc(din_27_ab0_1sc), .a1b1_1sc(din_27_ab1_1sc), .a1b2_1sc(din_27_ab2_1sc),
           .msk_a1b0(din_27_msk_ab0), .msk_a1b1(din_27_msk_ab1), .msk_a1b2(din_27_msk_ab2),
           .msk_a1b0_1sc(din_27_msk_ab0_1sc), .msk_a1b1_1sc(din_27_msk_ab1_1sc), .msk_a1b2_1sc(din_27_msk_ab2_1sc),

           .a2b0(din_29_ab0), .a2b1(din_29_ab1),
           .a2b0_1sc(din_29_ab0_1sc), .a2b1_1sc(din_29_ab1_1sc),
           .msk_a2b0(din_29_msk_ab0), .msk_a2b1(din_29_msk_ab1),
           .msk_a2b0_1sc(din_29_msk_ab0_1sc), .msk_a2b1_1sc(din_29_msk_ab1_1sc),
           
           .a3b0(din_31_ab0),
           .a3b0_1sc(din_31_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_26_calc (
           .clk(clk), .sign(din_signs_reg[26]), 
           .p(addr_6_26),
           .a0b0(din_26_ab0), .a0b1(din_26_ab1), .a0b2(din_26_ab2), .a0b3(din_26_ab3),
           .a0b0_1sc(din_26_ab0_1sc), .a0b1_1sc(din_26_ab1_1sc), .a0b2_1sc(din_26_ab2_1sc), .a0b3_1sc(din_26_ab3_1sc),
           .msk_a0b0(din_26_msk_ab0), .msk_a0b1(din_26_msk_ab1), .msk_a0b2(din_26_msk_ab2), .msk_a0b3(din_26_msk_ab3),
           .msk_a0b0_1sc(din_26_msk_ab0_1sc), .msk_a0b1_1sc(din_26_msk_ab1_1sc), .msk_a0b2_1sc(din_26_msk_ab2_1sc), .msk_a0b3_1sc(din_26_msk_ab3_1sc),

           .a1b0(din_28_ab0), .a1b1(din_28_ab1), .a1b2(din_28_ab2),
           .a1b0_1sc(din_28_ab0_1sc), .a1b1_1sc(din_28_ab1_1sc), .a1b2_1sc(din_28_ab2_1sc),
           .msk_a1b0(din_28_msk_ab0), .msk_a1b1(din_28_msk_ab1), .msk_a1b2(din_28_msk_ab2),
           .msk_a1b0_1sc(din_28_msk_ab0_1sc), .msk_a1b1_1sc(din_28_msk_ab1_1sc), .msk_a1b2_1sc(din_28_msk_ab2_1sc),

           .a2b0(din_30_ab0), .a2b1(din_30_ab1),
           .a2b0_1sc(din_30_ab0_1sc), .a2b1_1sc(din_30_ab1_1sc),
           .msk_a2b0(din_30_msk_ab0), .msk_a2b1(din_30_msk_ab1),
           .msk_a2b0_1sc(din_30_msk_ab0_1sc), .msk_a2b1_1sc(din_30_msk_ab1_1sc),
           
           .a3b0(din_32_ab0),
           .a3b0_1sc(din_32_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_27_calc (
           .clk(clk), .sign(din_signs_reg[27]), 
           .p(addr_6_27),
           .a0b0(din_27_ab0), .a0b1(din_27_ab1), .a0b2(din_27_ab2), .a0b3(din_27_ab3),
           .a0b0_1sc(din_27_ab0_1sc), .a0b1_1sc(din_27_ab1_1sc), .a0b2_1sc(din_27_ab2_1sc), .a0b3_1sc(din_27_ab3_1sc),
           .msk_a0b0(din_27_msk_ab0), .msk_a0b1(din_27_msk_ab1), .msk_a0b2(din_27_msk_ab2), .msk_a0b3(din_27_msk_ab3),
           .msk_a0b0_1sc(din_27_msk_ab0_1sc), .msk_a0b1_1sc(din_27_msk_ab1_1sc), .msk_a0b2_1sc(din_27_msk_ab2_1sc), .msk_a0b3_1sc(din_27_msk_ab3_1sc),

           .a1b0(din_29_ab0), .a1b1(din_29_ab1), .a1b2(din_29_ab2),
           .a1b0_1sc(din_29_ab0_1sc), .a1b1_1sc(din_29_ab1_1sc), .a1b2_1sc(din_29_ab2_1sc),
           .msk_a1b0(din_29_msk_ab0), .msk_a1b1(din_29_msk_ab1), .msk_a1b2(din_29_msk_ab2),
           .msk_a1b0_1sc(din_29_msk_ab0_1sc), .msk_a1b1_1sc(din_29_msk_ab1_1sc), .msk_a1b2_1sc(din_29_msk_ab2_1sc),

           .a2b0(din_31_ab0), .a2b1(din_31_ab1),
           .a2b0_1sc(din_31_ab0_1sc), .a2b1_1sc(din_31_ab1_1sc),
           .msk_a2b0(din_31_msk_ab0), .msk_a2b1(din_31_msk_ab1),
           .msk_a2b0_1sc(din_31_msk_ab0_1sc), .msk_a2b1_1sc(din_31_msk_ab1_1sc),
           
           .a3b0(din_33_ab0),
           .a3b0_1sc(din_33_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_28_calc (
           .clk(clk), .sign(din_signs_reg[28]), 
           .p(addr_6_28),
           .a0b0(din_28_ab0), .a0b1(din_28_ab1), .a0b2(din_28_ab2), .a0b3(din_28_ab3),
           .a0b0_1sc(din_28_ab0_1sc), .a0b1_1sc(din_28_ab1_1sc), .a0b2_1sc(din_28_ab2_1sc), .a0b3_1sc(din_28_ab3_1sc),
           .msk_a0b0(din_28_msk_ab0), .msk_a0b1(din_28_msk_ab1), .msk_a0b2(din_28_msk_ab2), .msk_a0b3(din_28_msk_ab3),
           .msk_a0b0_1sc(din_28_msk_ab0_1sc), .msk_a0b1_1sc(din_28_msk_ab1_1sc), .msk_a0b2_1sc(din_28_msk_ab2_1sc), .msk_a0b3_1sc(din_28_msk_ab3_1sc),

           .a1b0(din_30_ab0), .a1b1(din_30_ab1), .a1b2(din_30_ab2),
           .a1b0_1sc(din_30_ab0_1sc), .a1b1_1sc(din_30_ab1_1sc), .a1b2_1sc(din_30_ab2_1sc),
           .msk_a1b0(din_30_msk_ab0), .msk_a1b1(din_30_msk_ab1), .msk_a1b2(din_30_msk_ab2),
           .msk_a1b0_1sc(din_30_msk_ab0_1sc), .msk_a1b1_1sc(din_30_msk_ab1_1sc), .msk_a1b2_1sc(din_30_msk_ab2_1sc),

           .a2b0(din_32_ab0), .a2b1(din_32_ab1),
           .a2b0_1sc(din_32_ab0_1sc), .a2b1_1sc(din_32_ab1_1sc),
           .msk_a2b0(din_32_msk_ab0), .msk_a2b1(din_32_msk_ab1),
           .msk_a2b0_1sc(din_32_msk_ab0_1sc), .msk_a2b1_1sc(din_32_msk_ab1_1sc),
           
           .a3b0(din_34_ab0),
           .a3b0_1sc(din_34_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_29_calc (
           .clk(clk), .sign(din_signs_reg[29]), 
           .p(addr_6_29),
           .a0b0(din_29_ab0), .a0b1(din_29_ab1), .a0b2(din_29_ab2), .a0b3(din_29_ab3),
           .a0b0_1sc(din_29_ab0_1sc), .a0b1_1sc(din_29_ab1_1sc), .a0b2_1sc(din_29_ab2_1sc), .a0b3_1sc(din_29_ab3_1sc),
           .msk_a0b0(din_29_msk_ab0), .msk_a0b1(din_29_msk_ab1), .msk_a0b2(din_29_msk_ab2), .msk_a0b3(din_29_msk_ab3),
           .msk_a0b0_1sc(din_29_msk_ab0_1sc), .msk_a0b1_1sc(din_29_msk_ab1_1sc), .msk_a0b2_1sc(din_29_msk_ab2_1sc), .msk_a0b3_1sc(din_29_msk_ab3_1sc),

           .a1b0(din_31_ab0), .a1b1(din_31_ab1), .a1b2(din_31_ab2),
           .a1b0_1sc(din_31_ab0_1sc), .a1b1_1sc(din_31_ab1_1sc), .a1b2_1sc(din_31_ab2_1sc),
           .msk_a1b0(din_31_msk_ab0), .msk_a1b1(din_31_msk_ab1), .msk_a1b2(din_31_msk_ab2),
           .msk_a1b0_1sc(din_31_msk_ab0_1sc), .msk_a1b1_1sc(din_31_msk_ab1_1sc), .msk_a1b2_1sc(din_31_msk_ab2_1sc),

           .a2b0(din_33_ab0), .a2b1(din_33_ab1),
           .a2b0_1sc(din_33_ab0_1sc), .a2b1_1sc(din_33_ab1_1sc),
           .msk_a2b0(din_33_msk_ab0), .msk_a2b1(din_33_msk_ab1),
           .msk_a2b0_1sc(din_33_msk_ab0_1sc), .msk_a2b1_1sc(din_33_msk_ab1_1sc),
           
           .a3b0(din_35_ab0),
           .a3b0_1sc(din_35_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_30_calc (
           .clk(clk), .sign(din_signs_reg[30]), 
           .p(addr_6_30),
           .a0b0(din_30_ab0), .a0b1(din_30_ab1), .a0b2(din_30_ab2), .a0b3(din_30_ab3),
           .a0b0_1sc(din_30_ab0_1sc), .a0b1_1sc(din_30_ab1_1sc), .a0b2_1sc(din_30_ab2_1sc), .a0b3_1sc(din_30_ab3_1sc),
           .msk_a0b0(din_30_msk_ab0), .msk_a0b1(din_30_msk_ab1), .msk_a0b2(din_30_msk_ab2), .msk_a0b3(din_30_msk_ab3),
           .msk_a0b0_1sc(din_30_msk_ab0_1sc), .msk_a0b1_1sc(din_30_msk_ab1_1sc), .msk_a0b2_1sc(din_30_msk_ab2_1sc), .msk_a0b3_1sc(din_30_msk_ab3_1sc),

           .a1b0(din_32_ab0), .a1b1(din_32_ab1), .a1b2(din_32_ab2),
           .a1b0_1sc(din_32_ab0_1sc), .a1b1_1sc(din_32_ab1_1sc), .a1b2_1sc(din_32_ab2_1sc),
           .msk_a1b0(din_32_msk_ab0), .msk_a1b1(din_32_msk_ab1), .msk_a1b2(din_32_msk_ab2),
           .msk_a1b0_1sc(din_32_msk_ab0_1sc), .msk_a1b1_1sc(din_32_msk_ab1_1sc), .msk_a1b2_1sc(din_32_msk_ab2_1sc),

           .a2b0(din_34_ab0), .a2b1(din_34_ab1),
           .a2b0_1sc(din_34_ab0_1sc), .a2b1_1sc(din_34_ab1_1sc),
           .msk_a2b0(din_34_msk_ab0), .msk_a2b1(din_34_msk_ab1),
           .msk_a2b0_1sc(din_34_msk_ab0_1sc), .msk_a2b1_1sc(din_34_msk_ab1_1sc),
           
           .a3b0(din_36_ab0),
           .a3b0_1sc(din_36_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10)
) addr_6_31_calc (
           .clk(clk), .sign(din_signs_reg[31]), 
           .p(addr_6_31),
           .a0b0(din_31_ab0), .a0b1(din_31_ab1), .a0b2(din_31_ab2), .a0b3(din_31_ab3),
           .a0b0_1sc(din_31_ab0_1sc), .a0b1_1sc(din_31_ab1_1sc), .a0b2_1sc(din_31_ab2_1sc), .a0b3_1sc(din_31_ab3_1sc),
           .msk_a0b0(din_31_msk_ab0), .msk_a0b1(din_31_msk_ab1), .msk_a0b2(din_31_msk_ab2), .msk_a0b3(din_31_msk_ab3),
           .msk_a0b0_1sc(din_31_msk_ab0_1sc), .msk_a0b1_1sc(din_31_msk_ab1_1sc), .msk_a0b2_1sc(din_31_msk_ab2_1sc), .msk_a0b3_1sc(din_31_msk_ab3_1sc),

           .a1b0(din_33_ab0), .a1b1(din_33_ab1), .a1b2(din_33_ab2),
           .a1b0_1sc(din_33_ab0_1sc), .a1b1_1sc(din_33_ab1_1sc), .a1b2_1sc(din_33_ab2_1sc),
           .msk_a1b0(din_33_msk_ab0), .msk_a1b1(din_33_msk_ab1), .msk_a1b2(din_33_msk_ab2),
           .msk_a1b0_1sc(din_33_msk_ab0_1sc), .msk_a1b1_1sc(din_33_msk_ab1_1sc), .msk_a1b2_1sc(din_33_msk_ab2_1sc),

           .a2b0(din_35_ab0), .a2b1(din_35_ab1),
           .a2b0_1sc(din_35_ab0_1sc), .a2b1_1sc(din_35_ab1_1sc),
           .msk_a2b0(din_35_msk_ab0), .msk_a2b1(din_35_msk_ab1),
           .msk_a2b0_1sc(din_35_msk_ab0_1sc), .msk_a2b1_1sc(din_35_msk_ab1_1sc),
           
           .a3b0(din_37_ab0),
           .a3b0_1sc(din_37_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_0_calc (
           .clk(clk), .sign(din_signs_reg[0]), 
           .p(addr_7_0),
           .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
           .a0b0_1sc(din_0_ab0_1sc), .a0b1_1sc(din_0_ab1_1sc), .a0b2_1sc(din_0_ab2_1sc), .a0b3_1sc(din_0_ab3_1sc),
           .msk_a0b0(din_0_msk_ab0), .msk_a0b1(din_0_msk_ab1), .msk_a0b2(din_0_msk_ab2), .msk_a0b3(din_0_msk_ab3),
           .msk_a0b0_1sc(din_0_msk_ab0_1sc), .msk_a0b1_1sc(din_0_msk_ab1_1sc), .msk_a0b2_1sc(din_0_msk_ab2_1sc), .msk_a0b3_1sc(din_0_msk_ab3_1sc),

           .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2),
           .a1b0_1sc(din_2_ab0_1sc), .a1b1_1sc(din_2_ab1_1sc), .a1b2_1sc(din_2_ab2_1sc),
           .msk_a1b0(din_2_msk_ab0), .msk_a1b1(din_2_msk_ab1), .msk_a1b2(din_2_msk_ab2),
           .msk_a1b0_1sc(din_2_msk_ab0_1sc), .msk_a1b1_1sc(din_2_msk_ab1_1sc), .msk_a1b2_1sc(din_2_msk_ab2_1sc),

           .a2b0(din_4_ab0), .a2b1(din_4_ab1),
           .a2b0_1sc(din_4_ab0_1sc), .a2b1_1sc(din_4_ab1_1sc),
           .msk_a2b0(din_4_msk_ab0), .msk_a2b1(din_4_msk_ab1),
           .msk_a2b0_1sc(din_4_msk_ab0_1sc), .msk_a2b1_1sc(din_4_msk_ab1_1sc),
           
           .a3b0(din_6_ab0),
           .a3b0_1sc(din_6_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_1_calc (
           .clk(clk), .sign(din_signs_reg[1]), 
           .p(addr_7_1),
           .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
           .a0b0_1sc(din_1_ab0_1sc), .a0b1_1sc(din_1_ab1_1sc), .a0b2_1sc(din_1_ab2_1sc), .a0b3_1sc(din_1_ab3_1sc),
           .msk_a0b0(din_1_msk_ab0), .msk_a0b1(din_1_msk_ab1), .msk_a0b2(din_1_msk_ab2), .msk_a0b3(din_1_msk_ab3),
           .msk_a0b0_1sc(din_1_msk_ab0_1sc), .msk_a0b1_1sc(din_1_msk_ab1_1sc), .msk_a0b2_1sc(din_1_msk_ab2_1sc), .msk_a0b3_1sc(din_1_msk_ab3_1sc),

           .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2),
           .a1b0_1sc(din_3_ab0_1sc), .a1b1_1sc(din_3_ab1_1sc), .a1b2_1sc(din_3_ab2_1sc),
           .msk_a1b0(din_3_msk_ab0), .msk_a1b1(din_3_msk_ab1), .msk_a1b2(din_3_msk_ab2),
           .msk_a1b0_1sc(din_3_msk_ab0_1sc), .msk_a1b1_1sc(din_3_msk_ab1_1sc), .msk_a1b2_1sc(din_3_msk_ab2_1sc),

           .a2b0(din_5_ab0), .a2b1(din_5_ab1),
           .a2b0_1sc(din_5_ab0_1sc), .a2b1_1sc(din_5_ab1_1sc),
           .msk_a2b0(din_5_msk_ab0), .msk_a2b1(din_5_msk_ab1),
           .msk_a2b0_1sc(din_5_msk_ab0_1sc), .msk_a2b1_1sc(din_5_msk_ab1_1sc),
           
           .a3b0(din_7_ab0),
           .a3b0_1sc(din_7_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_2_calc (
           .clk(clk), .sign(din_signs_reg[2]), 
           .p(addr_7_2),
           .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
           .a0b0_1sc(din_2_ab0_1sc), .a0b1_1sc(din_2_ab1_1sc), .a0b2_1sc(din_2_ab2_1sc), .a0b3_1sc(din_2_ab3_1sc),
           .msk_a0b0(din_2_msk_ab0), .msk_a0b1(din_2_msk_ab1), .msk_a0b2(din_2_msk_ab2), .msk_a0b3(din_2_msk_ab3),
           .msk_a0b0_1sc(din_2_msk_ab0_1sc), .msk_a0b1_1sc(din_2_msk_ab1_1sc), .msk_a0b2_1sc(din_2_msk_ab2_1sc), .msk_a0b3_1sc(din_2_msk_ab3_1sc),

           .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2),
           .a1b0_1sc(din_4_ab0_1sc), .a1b1_1sc(din_4_ab1_1sc), .a1b2_1sc(din_4_ab2_1sc),
           .msk_a1b0(din_4_msk_ab0), .msk_a1b1(din_4_msk_ab1), .msk_a1b2(din_4_msk_ab2),
           .msk_a1b0_1sc(din_4_msk_ab0_1sc), .msk_a1b1_1sc(din_4_msk_ab1_1sc), .msk_a1b2_1sc(din_4_msk_ab2_1sc),

           .a2b0(din_6_ab0), .a2b1(din_6_ab1),
           .a2b0_1sc(din_6_ab0_1sc), .a2b1_1sc(din_6_ab1_1sc),
           .msk_a2b0(din_6_msk_ab0), .msk_a2b1(din_6_msk_ab1),
           .msk_a2b0_1sc(din_6_msk_ab0_1sc), .msk_a2b1_1sc(din_6_msk_ab1_1sc),
           
           .a3b0(din_8_ab0),
           .a3b0_1sc(din_8_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_3_calc (
           .clk(clk), .sign(din_signs_reg[3]), 
           .p(addr_7_3),
           .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
           .a0b0_1sc(din_3_ab0_1sc), .a0b1_1sc(din_3_ab1_1sc), .a0b2_1sc(din_3_ab2_1sc), .a0b3_1sc(din_3_ab3_1sc),
           .msk_a0b0(din_3_msk_ab0), .msk_a0b1(din_3_msk_ab1), .msk_a0b2(din_3_msk_ab2), .msk_a0b3(din_3_msk_ab3),
           .msk_a0b0_1sc(din_3_msk_ab0_1sc), .msk_a0b1_1sc(din_3_msk_ab1_1sc), .msk_a0b2_1sc(din_3_msk_ab2_1sc), .msk_a0b3_1sc(din_3_msk_ab3_1sc),

           .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2),
           .a1b0_1sc(din_5_ab0_1sc), .a1b1_1sc(din_5_ab1_1sc), .a1b2_1sc(din_5_ab2_1sc),
           .msk_a1b0(din_5_msk_ab0), .msk_a1b1(din_5_msk_ab1), .msk_a1b2(din_5_msk_ab2),
           .msk_a1b0_1sc(din_5_msk_ab0_1sc), .msk_a1b1_1sc(din_5_msk_ab1_1sc), .msk_a1b2_1sc(din_5_msk_ab2_1sc),

           .a2b0(din_7_ab0), .a2b1(din_7_ab1),
           .a2b0_1sc(din_7_ab0_1sc), .a2b1_1sc(din_7_ab1_1sc),
           .msk_a2b0(din_7_msk_ab0), .msk_a2b1(din_7_msk_ab1),
           .msk_a2b0_1sc(din_7_msk_ab0_1sc), .msk_a2b1_1sc(din_7_msk_ab1_1sc),
           
           .a3b0(din_9_ab0),
           .a3b0_1sc(din_9_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_4_calc (
           .clk(clk), .sign(din_signs_reg[4]), 
           .p(addr_7_4),
           .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
           .a0b0_1sc(din_4_ab0_1sc), .a0b1_1sc(din_4_ab1_1sc), .a0b2_1sc(din_4_ab2_1sc), .a0b3_1sc(din_4_ab3_1sc),
           .msk_a0b0(din_4_msk_ab0), .msk_a0b1(din_4_msk_ab1), .msk_a0b2(din_4_msk_ab2), .msk_a0b3(din_4_msk_ab3),
           .msk_a0b0_1sc(din_4_msk_ab0_1sc), .msk_a0b1_1sc(din_4_msk_ab1_1sc), .msk_a0b2_1sc(din_4_msk_ab2_1sc), .msk_a0b3_1sc(din_4_msk_ab3_1sc),

           .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2),
           .a1b0_1sc(din_6_ab0_1sc), .a1b1_1sc(din_6_ab1_1sc), .a1b2_1sc(din_6_ab2_1sc),
           .msk_a1b0(din_6_msk_ab0), .msk_a1b1(din_6_msk_ab1), .msk_a1b2(din_6_msk_ab2),
           .msk_a1b0_1sc(din_6_msk_ab0_1sc), .msk_a1b1_1sc(din_6_msk_ab1_1sc), .msk_a1b2_1sc(din_6_msk_ab2_1sc),

           .a2b0(din_8_ab0), .a2b1(din_8_ab1),
           .a2b0_1sc(din_8_ab0_1sc), .a2b1_1sc(din_8_ab1_1sc),
           .msk_a2b0(din_8_msk_ab0), .msk_a2b1(din_8_msk_ab1),
           .msk_a2b0_1sc(din_8_msk_ab0_1sc), .msk_a2b1_1sc(din_8_msk_ab1_1sc),
           
           .a3b0(din_10_ab0),
           .a3b0_1sc(din_10_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_5_calc (
           .clk(clk), .sign(din_signs_reg[5]), 
           .p(addr_7_5),
           .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
           .a0b0_1sc(din_5_ab0_1sc), .a0b1_1sc(din_5_ab1_1sc), .a0b2_1sc(din_5_ab2_1sc), .a0b3_1sc(din_5_ab3_1sc),
           .msk_a0b0(din_5_msk_ab0), .msk_a0b1(din_5_msk_ab1), .msk_a0b2(din_5_msk_ab2), .msk_a0b3(din_5_msk_ab3),
           .msk_a0b0_1sc(din_5_msk_ab0_1sc), .msk_a0b1_1sc(din_5_msk_ab1_1sc), .msk_a0b2_1sc(din_5_msk_ab2_1sc), .msk_a0b3_1sc(din_5_msk_ab3_1sc),

           .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2),
           .a1b0_1sc(din_7_ab0_1sc), .a1b1_1sc(din_7_ab1_1sc), .a1b2_1sc(din_7_ab2_1sc),
           .msk_a1b0(din_7_msk_ab0), .msk_a1b1(din_7_msk_ab1), .msk_a1b2(din_7_msk_ab2),
           .msk_a1b0_1sc(din_7_msk_ab0_1sc), .msk_a1b1_1sc(din_7_msk_ab1_1sc), .msk_a1b2_1sc(din_7_msk_ab2_1sc),

           .a2b0(din_9_ab0), .a2b1(din_9_ab1),
           .a2b0_1sc(din_9_ab0_1sc), .a2b1_1sc(din_9_ab1_1sc),
           .msk_a2b0(din_9_msk_ab0), .msk_a2b1(din_9_msk_ab1),
           .msk_a2b0_1sc(din_9_msk_ab0_1sc), .msk_a2b1_1sc(din_9_msk_ab1_1sc),
           
           .a3b0(din_11_ab0),
           .a3b0_1sc(din_11_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_6_calc (
           .clk(clk), .sign(din_signs_reg[6]), 
           .p(addr_7_6),
           .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
           .a0b0_1sc(din_6_ab0_1sc), .a0b1_1sc(din_6_ab1_1sc), .a0b2_1sc(din_6_ab2_1sc), .a0b3_1sc(din_6_ab3_1sc),
           .msk_a0b0(din_6_msk_ab0), .msk_a0b1(din_6_msk_ab1), .msk_a0b2(din_6_msk_ab2), .msk_a0b3(din_6_msk_ab3),
           .msk_a0b0_1sc(din_6_msk_ab0_1sc), .msk_a0b1_1sc(din_6_msk_ab1_1sc), .msk_a0b2_1sc(din_6_msk_ab2_1sc), .msk_a0b3_1sc(din_6_msk_ab3_1sc),

           .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2),
           .a1b0_1sc(din_8_ab0_1sc), .a1b1_1sc(din_8_ab1_1sc), .a1b2_1sc(din_8_ab2_1sc),
           .msk_a1b0(din_8_msk_ab0), .msk_a1b1(din_8_msk_ab1), .msk_a1b2(din_8_msk_ab2),
           .msk_a1b0_1sc(din_8_msk_ab0_1sc), .msk_a1b1_1sc(din_8_msk_ab1_1sc), .msk_a1b2_1sc(din_8_msk_ab2_1sc),

           .a2b0(din_10_ab0), .a2b1(din_10_ab1),
           .a2b0_1sc(din_10_ab0_1sc), .a2b1_1sc(din_10_ab1_1sc),
           .msk_a2b0(din_10_msk_ab0), .msk_a2b1(din_10_msk_ab1),
           .msk_a2b0_1sc(din_10_msk_ab0_1sc), .msk_a2b1_1sc(din_10_msk_ab1_1sc),
           
           .a3b0(din_12_ab0),
           .a3b0_1sc(din_12_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_7_calc (
           .clk(clk), .sign(din_signs_reg[7]), 
           .p(addr_7_7),
           .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
           .a0b0_1sc(din_7_ab0_1sc), .a0b1_1sc(din_7_ab1_1sc), .a0b2_1sc(din_7_ab2_1sc), .a0b3_1sc(din_7_ab3_1sc),
           .msk_a0b0(din_7_msk_ab0), .msk_a0b1(din_7_msk_ab1), .msk_a0b2(din_7_msk_ab2), .msk_a0b3(din_7_msk_ab3),
           .msk_a0b0_1sc(din_7_msk_ab0_1sc), .msk_a0b1_1sc(din_7_msk_ab1_1sc), .msk_a0b2_1sc(din_7_msk_ab2_1sc), .msk_a0b3_1sc(din_7_msk_ab3_1sc),

           .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2),
           .a1b0_1sc(din_9_ab0_1sc), .a1b1_1sc(din_9_ab1_1sc), .a1b2_1sc(din_9_ab2_1sc),
           .msk_a1b0(din_9_msk_ab0), .msk_a1b1(din_9_msk_ab1), .msk_a1b2(din_9_msk_ab2),
           .msk_a1b0_1sc(din_9_msk_ab0_1sc), .msk_a1b1_1sc(din_9_msk_ab1_1sc), .msk_a1b2_1sc(din_9_msk_ab2_1sc),

           .a2b0(din_11_ab0), .a2b1(din_11_ab1),
           .a2b0_1sc(din_11_ab0_1sc), .a2b1_1sc(din_11_ab1_1sc),
           .msk_a2b0(din_11_msk_ab0), .msk_a2b1(din_11_msk_ab1),
           .msk_a2b0_1sc(din_11_msk_ab0_1sc), .msk_a2b1_1sc(din_11_msk_ab1_1sc),
           
           .a3b0(din_13_ab0),
           .a3b0_1sc(din_13_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_8_calc (
           .clk(clk), .sign(din_signs_reg[8]), 
           .p(addr_7_8),
           .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
           .a0b0_1sc(din_8_ab0_1sc), .a0b1_1sc(din_8_ab1_1sc), .a0b2_1sc(din_8_ab2_1sc), .a0b3_1sc(din_8_ab3_1sc),
           .msk_a0b0(din_8_msk_ab0), .msk_a0b1(din_8_msk_ab1), .msk_a0b2(din_8_msk_ab2), .msk_a0b3(din_8_msk_ab3),
           .msk_a0b0_1sc(din_8_msk_ab0_1sc), .msk_a0b1_1sc(din_8_msk_ab1_1sc), .msk_a0b2_1sc(din_8_msk_ab2_1sc), .msk_a0b3_1sc(din_8_msk_ab3_1sc),

           .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2),
           .a1b0_1sc(din_10_ab0_1sc), .a1b1_1sc(din_10_ab1_1sc), .a1b2_1sc(din_10_ab2_1sc),
           .msk_a1b0(din_10_msk_ab0), .msk_a1b1(din_10_msk_ab1), .msk_a1b2(din_10_msk_ab2),
           .msk_a1b0_1sc(din_10_msk_ab0_1sc), .msk_a1b1_1sc(din_10_msk_ab1_1sc), .msk_a1b2_1sc(din_10_msk_ab2_1sc),

           .a2b0(din_12_ab0), .a2b1(din_12_ab1),
           .a2b0_1sc(din_12_ab0_1sc), .a2b1_1sc(din_12_ab1_1sc),
           .msk_a2b0(din_12_msk_ab0), .msk_a2b1(din_12_msk_ab1),
           .msk_a2b0_1sc(din_12_msk_ab0_1sc), .msk_a2b1_1sc(din_12_msk_ab1_1sc),
           
           .a3b0(din_14_ab0),
           .a3b0_1sc(din_14_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_9_calc (
           .clk(clk), .sign(din_signs_reg[9]), 
           .p(addr_7_9),
           .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
           .a0b0_1sc(din_9_ab0_1sc), .a0b1_1sc(din_9_ab1_1sc), .a0b2_1sc(din_9_ab2_1sc), .a0b3_1sc(din_9_ab3_1sc),
           .msk_a0b0(din_9_msk_ab0), .msk_a0b1(din_9_msk_ab1), .msk_a0b2(din_9_msk_ab2), .msk_a0b3(din_9_msk_ab3),
           .msk_a0b0_1sc(din_9_msk_ab0_1sc), .msk_a0b1_1sc(din_9_msk_ab1_1sc), .msk_a0b2_1sc(din_9_msk_ab2_1sc), .msk_a0b3_1sc(din_9_msk_ab3_1sc),

           .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2),
           .a1b0_1sc(din_11_ab0_1sc), .a1b1_1sc(din_11_ab1_1sc), .a1b2_1sc(din_11_ab2_1sc),
           .msk_a1b0(din_11_msk_ab0), .msk_a1b1(din_11_msk_ab1), .msk_a1b2(din_11_msk_ab2),
           .msk_a1b0_1sc(din_11_msk_ab0_1sc), .msk_a1b1_1sc(din_11_msk_ab1_1sc), .msk_a1b2_1sc(din_11_msk_ab2_1sc),

           .a2b0(din_13_ab0), .a2b1(din_13_ab1),
           .a2b0_1sc(din_13_ab0_1sc), .a2b1_1sc(din_13_ab1_1sc),
           .msk_a2b0(din_13_msk_ab0), .msk_a2b1(din_13_msk_ab1),
           .msk_a2b0_1sc(din_13_msk_ab0_1sc), .msk_a2b1_1sc(din_13_msk_ab1_1sc),
           
           .a3b0(din_15_ab0),
           .a3b0_1sc(din_15_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_10_calc (
           .clk(clk), .sign(din_signs_reg[10]), 
           .p(addr_7_10),
           .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
           .a0b0_1sc(din_10_ab0_1sc), .a0b1_1sc(din_10_ab1_1sc), .a0b2_1sc(din_10_ab2_1sc), .a0b3_1sc(din_10_ab3_1sc),
           .msk_a0b0(din_10_msk_ab0), .msk_a0b1(din_10_msk_ab1), .msk_a0b2(din_10_msk_ab2), .msk_a0b3(din_10_msk_ab3),
           .msk_a0b0_1sc(din_10_msk_ab0_1sc), .msk_a0b1_1sc(din_10_msk_ab1_1sc), .msk_a0b2_1sc(din_10_msk_ab2_1sc), .msk_a0b3_1sc(din_10_msk_ab3_1sc),

           .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2),
           .a1b0_1sc(din_12_ab0_1sc), .a1b1_1sc(din_12_ab1_1sc), .a1b2_1sc(din_12_ab2_1sc),
           .msk_a1b0(din_12_msk_ab0), .msk_a1b1(din_12_msk_ab1), .msk_a1b2(din_12_msk_ab2),
           .msk_a1b0_1sc(din_12_msk_ab0_1sc), .msk_a1b1_1sc(din_12_msk_ab1_1sc), .msk_a1b2_1sc(din_12_msk_ab2_1sc),

           .a2b0(din_14_ab0), .a2b1(din_14_ab1),
           .a2b0_1sc(din_14_ab0_1sc), .a2b1_1sc(din_14_ab1_1sc),
           .msk_a2b0(din_14_msk_ab0), .msk_a2b1(din_14_msk_ab1),
           .msk_a2b0_1sc(din_14_msk_ab0_1sc), .msk_a2b1_1sc(din_14_msk_ab1_1sc),
           
           .a3b0(din_16_ab0),
           .a3b0_1sc(din_16_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_11_calc (
           .clk(clk), .sign(din_signs_reg[11]), 
           .p(addr_7_11),
           .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
           .a0b0_1sc(din_11_ab0_1sc), .a0b1_1sc(din_11_ab1_1sc), .a0b2_1sc(din_11_ab2_1sc), .a0b3_1sc(din_11_ab3_1sc),
           .msk_a0b0(din_11_msk_ab0), .msk_a0b1(din_11_msk_ab1), .msk_a0b2(din_11_msk_ab2), .msk_a0b3(din_11_msk_ab3),
           .msk_a0b0_1sc(din_11_msk_ab0_1sc), .msk_a0b1_1sc(din_11_msk_ab1_1sc), .msk_a0b2_1sc(din_11_msk_ab2_1sc), .msk_a0b3_1sc(din_11_msk_ab3_1sc),

           .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2),
           .a1b0_1sc(din_13_ab0_1sc), .a1b1_1sc(din_13_ab1_1sc), .a1b2_1sc(din_13_ab2_1sc),
           .msk_a1b0(din_13_msk_ab0), .msk_a1b1(din_13_msk_ab1), .msk_a1b2(din_13_msk_ab2),
           .msk_a1b0_1sc(din_13_msk_ab0_1sc), .msk_a1b1_1sc(din_13_msk_ab1_1sc), .msk_a1b2_1sc(din_13_msk_ab2_1sc),

           .a2b0(din_15_ab0), .a2b1(din_15_ab1),
           .a2b0_1sc(din_15_ab0_1sc), .a2b1_1sc(din_15_ab1_1sc),
           .msk_a2b0(din_15_msk_ab0), .msk_a2b1(din_15_msk_ab1),
           .msk_a2b0_1sc(din_15_msk_ab0_1sc), .msk_a2b1_1sc(din_15_msk_ab1_1sc),
           
           .a3b0(din_17_ab0),
           .a3b0_1sc(din_17_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_12_calc (
           .clk(clk), .sign(din_signs_reg[12]), 
           .p(addr_7_12),
           .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
           .a0b0_1sc(din_12_ab0_1sc), .a0b1_1sc(din_12_ab1_1sc), .a0b2_1sc(din_12_ab2_1sc), .a0b3_1sc(din_12_ab3_1sc),
           .msk_a0b0(din_12_msk_ab0), .msk_a0b1(din_12_msk_ab1), .msk_a0b2(din_12_msk_ab2), .msk_a0b3(din_12_msk_ab3),
           .msk_a0b0_1sc(din_12_msk_ab0_1sc), .msk_a0b1_1sc(din_12_msk_ab1_1sc), .msk_a0b2_1sc(din_12_msk_ab2_1sc), .msk_a0b3_1sc(din_12_msk_ab3_1sc),

           .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2),
           .a1b0_1sc(din_14_ab0_1sc), .a1b1_1sc(din_14_ab1_1sc), .a1b2_1sc(din_14_ab2_1sc),
           .msk_a1b0(din_14_msk_ab0), .msk_a1b1(din_14_msk_ab1), .msk_a1b2(din_14_msk_ab2),
           .msk_a1b0_1sc(din_14_msk_ab0_1sc), .msk_a1b1_1sc(din_14_msk_ab1_1sc), .msk_a1b2_1sc(din_14_msk_ab2_1sc),

           .a2b0(din_16_ab0), .a2b1(din_16_ab1),
           .a2b0_1sc(din_16_ab0_1sc), .a2b1_1sc(din_16_ab1_1sc),
           .msk_a2b0(din_16_msk_ab0), .msk_a2b1(din_16_msk_ab1),
           .msk_a2b0_1sc(din_16_msk_ab0_1sc), .msk_a2b1_1sc(din_16_msk_ab1_1sc),
           
           .a3b0(din_18_ab0),
           .a3b0_1sc(din_18_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_13_calc (
           .clk(clk), .sign(din_signs_reg[13]), 
           .p(addr_7_13),
           .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
           .a0b0_1sc(din_13_ab0_1sc), .a0b1_1sc(din_13_ab1_1sc), .a0b2_1sc(din_13_ab2_1sc), .a0b3_1sc(din_13_ab3_1sc),
           .msk_a0b0(din_13_msk_ab0), .msk_a0b1(din_13_msk_ab1), .msk_a0b2(din_13_msk_ab2), .msk_a0b3(din_13_msk_ab3),
           .msk_a0b0_1sc(din_13_msk_ab0_1sc), .msk_a0b1_1sc(din_13_msk_ab1_1sc), .msk_a0b2_1sc(din_13_msk_ab2_1sc), .msk_a0b3_1sc(din_13_msk_ab3_1sc),

           .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2),
           .a1b0_1sc(din_15_ab0_1sc), .a1b1_1sc(din_15_ab1_1sc), .a1b2_1sc(din_15_ab2_1sc),
           .msk_a1b0(din_15_msk_ab0), .msk_a1b1(din_15_msk_ab1), .msk_a1b2(din_15_msk_ab2),
           .msk_a1b0_1sc(din_15_msk_ab0_1sc), .msk_a1b1_1sc(din_15_msk_ab1_1sc), .msk_a1b2_1sc(din_15_msk_ab2_1sc),

           .a2b0(din_17_ab0), .a2b1(din_17_ab1),
           .a2b0_1sc(din_17_ab0_1sc), .a2b1_1sc(din_17_ab1_1sc),
           .msk_a2b0(din_17_msk_ab0), .msk_a2b1(din_17_msk_ab1),
           .msk_a2b0_1sc(din_17_msk_ab0_1sc), .msk_a2b1_1sc(din_17_msk_ab1_1sc),
           
           .a3b0(din_19_ab0),
           .a3b0_1sc(din_19_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_14_calc (
           .clk(clk), .sign(din_signs_reg[14]), 
           .p(addr_7_14),
           .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
           .a0b0_1sc(din_14_ab0_1sc), .a0b1_1sc(din_14_ab1_1sc), .a0b2_1sc(din_14_ab2_1sc), .a0b3_1sc(din_14_ab3_1sc),
           .msk_a0b0(din_14_msk_ab0), .msk_a0b1(din_14_msk_ab1), .msk_a0b2(din_14_msk_ab2), .msk_a0b3(din_14_msk_ab3),
           .msk_a0b0_1sc(din_14_msk_ab0_1sc), .msk_a0b1_1sc(din_14_msk_ab1_1sc), .msk_a0b2_1sc(din_14_msk_ab2_1sc), .msk_a0b3_1sc(din_14_msk_ab3_1sc),

           .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2),
           .a1b0_1sc(din_16_ab0_1sc), .a1b1_1sc(din_16_ab1_1sc), .a1b2_1sc(din_16_ab2_1sc),
           .msk_a1b0(din_16_msk_ab0), .msk_a1b1(din_16_msk_ab1), .msk_a1b2(din_16_msk_ab2),
           .msk_a1b0_1sc(din_16_msk_ab0_1sc), .msk_a1b1_1sc(din_16_msk_ab1_1sc), .msk_a1b2_1sc(din_16_msk_ab2_1sc),

           .a2b0(din_18_ab0), .a2b1(din_18_ab1),
           .a2b0_1sc(din_18_ab0_1sc), .a2b1_1sc(din_18_ab1_1sc),
           .msk_a2b0(din_18_msk_ab0), .msk_a2b1(din_18_msk_ab1),
           .msk_a2b0_1sc(din_18_msk_ab0_1sc), .msk_a2b1_1sc(din_18_msk_ab1_1sc),
           
           .a3b0(din_20_ab0),
           .a3b0_1sc(din_20_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_15_calc (
           .clk(clk), .sign(din_signs_reg[15]), 
           .p(addr_7_15),
           .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
           .a0b0_1sc(din_15_ab0_1sc), .a0b1_1sc(din_15_ab1_1sc), .a0b2_1sc(din_15_ab2_1sc), .a0b3_1sc(din_15_ab3_1sc),
           .msk_a0b0(din_15_msk_ab0), .msk_a0b1(din_15_msk_ab1), .msk_a0b2(din_15_msk_ab2), .msk_a0b3(din_15_msk_ab3),
           .msk_a0b0_1sc(din_15_msk_ab0_1sc), .msk_a0b1_1sc(din_15_msk_ab1_1sc), .msk_a0b2_1sc(din_15_msk_ab2_1sc), .msk_a0b3_1sc(din_15_msk_ab3_1sc),

           .a1b0(din_17_ab0), .a1b1(din_17_ab1), .a1b2(din_17_ab2),
           .a1b0_1sc(din_17_ab0_1sc), .a1b1_1sc(din_17_ab1_1sc), .a1b2_1sc(din_17_ab2_1sc),
           .msk_a1b0(din_17_msk_ab0), .msk_a1b1(din_17_msk_ab1), .msk_a1b2(din_17_msk_ab2),
           .msk_a1b0_1sc(din_17_msk_ab0_1sc), .msk_a1b1_1sc(din_17_msk_ab1_1sc), .msk_a1b2_1sc(din_17_msk_ab2_1sc),

           .a2b0(din_19_ab0), .a2b1(din_19_ab1),
           .a2b0_1sc(din_19_ab0_1sc), .a2b1_1sc(din_19_ab1_1sc),
           .msk_a2b0(din_19_msk_ab0), .msk_a2b1(din_19_msk_ab1),
           .msk_a2b0_1sc(din_19_msk_ab0_1sc), .msk_a2b1_1sc(din_19_msk_ab1_1sc),
           
           .a3b0(din_21_ab0),
           .a3b0_1sc(din_21_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_16_calc (
           .clk(clk), .sign(din_signs_reg[16]), 
           .p(addr_7_16),
           .a0b0(din_16_ab0), .a0b1(din_16_ab1), .a0b2(din_16_ab2), .a0b3(din_16_ab3),
           .a0b0_1sc(din_16_ab0_1sc), .a0b1_1sc(din_16_ab1_1sc), .a0b2_1sc(din_16_ab2_1sc), .a0b3_1sc(din_16_ab3_1sc),
           .msk_a0b0(din_16_msk_ab0), .msk_a0b1(din_16_msk_ab1), .msk_a0b2(din_16_msk_ab2), .msk_a0b3(din_16_msk_ab3),
           .msk_a0b0_1sc(din_16_msk_ab0_1sc), .msk_a0b1_1sc(din_16_msk_ab1_1sc), .msk_a0b2_1sc(din_16_msk_ab2_1sc), .msk_a0b3_1sc(din_16_msk_ab3_1sc),

           .a1b0(din_18_ab0), .a1b1(din_18_ab1), .a1b2(din_18_ab2),
           .a1b0_1sc(din_18_ab0_1sc), .a1b1_1sc(din_18_ab1_1sc), .a1b2_1sc(din_18_ab2_1sc),
           .msk_a1b0(din_18_msk_ab0), .msk_a1b1(din_18_msk_ab1), .msk_a1b2(din_18_msk_ab2),
           .msk_a1b0_1sc(din_18_msk_ab0_1sc), .msk_a1b1_1sc(din_18_msk_ab1_1sc), .msk_a1b2_1sc(din_18_msk_ab2_1sc),

           .a2b0(din_20_ab0), .a2b1(din_20_ab1),
           .a2b0_1sc(din_20_ab0_1sc), .a2b1_1sc(din_20_ab1_1sc),
           .msk_a2b0(din_20_msk_ab0), .msk_a2b1(din_20_msk_ab1),
           .msk_a2b0_1sc(din_20_msk_ab0_1sc), .msk_a2b1_1sc(din_20_msk_ab1_1sc),
           
           .a3b0(din_22_ab0),
           .a3b0_1sc(din_22_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_17_calc (
           .clk(clk), .sign(din_signs_reg[17]), 
           .p(addr_7_17),
           .a0b0(din_17_ab0), .a0b1(din_17_ab1), .a0b2(din_17_ab2), .a0b3(din_17_ab3),
           .a0b0_1sc(din_17_ab0_1sc), .a0b1_1sc(din_17_ab1_1sc), .a0b2_1sc(din_17_ab2_1sc), .a0b3_1sc(din_17_ab3_1sc),
           .msk_a0b0(din_17_msk_ab0), .msk_a0b1(din_17_msk_ab1), .msk_a0b2(din_17_msk_ab2), .msk_a0b3(din_17_msk_ab3),
           .msk_a0b0_1sc(din_17_msk_ab0_1sc), .msk_a0b1_1sc(din_17_msk_ab1_1sc), .msk_a0b2_1sc(din_17_msk_ab2_1sc), .msk_a0b3_1sc(din_17_msk_ab3_1sc),

           .a1b0(din_19_ab0), .a1b1(din_19_ab1), .a1b2(din_19_ab2),
           .a1b0_1sc(din_19_ab0_1sc), .a1b1_1sc(din_19_ab1_1sc), .a1b2_1sc(din_19_ab2_1sc),
           .msk_a1b0(din_19_msk_ab0), .msk_a1b1(din_19_msk_ab1), .msk_a1b2(din_19_msk_ab2),
           .msk_a1b0_1sc(din_19_msk_ab0_1sc), .msk_a1b1_1sc(din_19_msk_ab1_1sc), .msk_a1b2_1sc(din_19_msk_ab2_1sc),

           .a2b0(din_21_ab0), .a2b1(din_21_ab1),
           .a2b0_1sc(din_21_ab0_1sc), .a2b1_1sc(din_21_ab1_1sc),
           .msk_a2b0(din_21_msk_ab0), .msk_a2b1(din_21_msk_ab1),
           .msk_a2b0_1sc(din_21_msk_ab0_1sc), .msk_a2b1_1sc(din_21_msk_ab1_1sc),
           
           .a3b0(din_23_ab0),
           .a3b0_1sc(din_23_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_18_calc (
           .clk(clk), .sign(din_signs_reg[18]), 
           .p(addr_7_18),
           .a0b0(din_18_ab0), .a0b1(din_18_ab1), .a0b2(din_18_ab2), .a0b3(din_18_ab3),
           .a0b0_1sc(din_18_ab0_1sc), .a0b1_1sc(din_18_ab1_1sc), .a0b2_1sc(din_18_ab2_1sc), .a0b3_1sc(din_18_ab3_1sc),
           .msk_a0b0(din_18_msk_ab0), .msk_a0b1(din_18_msk_ab1), .msk_a0b2(din_18_msk_ab2), .msk_a0b3(din_18_msk_ab3),
           .msk_a0b0_1sc(din_18_msk_ab0_1sc), .msk_a0b1_1sc(din_18_msk_ab1_1sc), .msk_a0b2_1sc(din_18_msk_ab2_1sc), .msk_a0b3_1sc(din_18_msk_ab3_1sc),

           .a1b0(din_20_ab0), .a1b1(din_20_ab1), .a1b2(din_20_ab2),
           .a1b0_1sc(din_20_ab0_1sc), .a1b1_1sc(din_20_ab1_1sc), .a1b2_1sc(din_20_ab2_1sc),
           .msk_a1b0(din_20_msk_ab0), .msk_a1b1(din_20_msk_ab1), .msk_a1b2(din_20_msk_ab2),
           .msk_a1b0_1sc(din_20_msk_ab0_1sc), .msk_a1b1_1sc(din_20_msk_ab1_1sc), .msk_a1b2_1sc(din_20_msk_ab2_1sc),

           .a2b0(din_22_ab0), .a2b1(din_22_ab1),
           .a2b0_1sc(din_22_ab0_1sc), .a2b1_1sc(din_22_ab1_1sc),
           .msk_a2b0(din_22_msk_ab0), .msk_a2b1(din_22_msk_ab1),
           .msk_a2b0_1sc(din_22_msk_ab0_1sc), .msk_a2b1_1sc(din_22_msk_ab1_1sc),
           
           .a3b0(din_24_ab0),
           .a3b0_1sc(din_24_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_19_calc (
           .clk(clk), .sign(din_signs_reg[19]), 
           .p(addr_7_19),
           .a0b0(din_19_ab0), .a0b1(din_19_ab1), .a0b2(din_19_ab2), .a0b3(din_19_ab3),
           .a0b0_1sc(din_19_ab0_1sc), .a0b1_1sc(din_19_ab1_1sc), .a0b2_1sc(din_19_ab2_1sc), .a0b3_1sc(din_19_ab3_1sc),
           .msk_a0b0(din_19_msk_ab0), .msk_a0b1(din_19_msk_ab1), .msk_a0b2(din_19_msk_ab2), .msk_a0b3(din_19_msk_ab3),
           .msk_a0b0_1sc(din_19_msk_ab0_1sc), .msk_a0b1_1sc(din_19_msk_ab1_1sc), .msk_a0b2_1sc(din_19_msk_ab2_1sc), .msk_a0b3_1sc(din_19_msk_ab3_1sc),

           .a1b0(din_21_ab0), .a1b1(din_21_ab1), .a1b2(din_21_ab2),
           .a1b0_1sc(din_21_ab0_1sc), .a1b1_1sc(din_21_ab1_1sc), .a1b2_1sc(din_21_ab2_1sc),
           .msk_a1b0(din_21_msk_ab0), .msk_a1b1(din_21_msk_ab1), .msk_a1b2(din_21_msk_ab2),
           .msk_a1b0_1sc(din_21_msk_ab0_1sc), .msk_a1b1_1sc(din_21_msk_ab1_1sc), .msk_a1b2_1sc(din_21_msk_ab2_1sc),

           .a2b0(din_23_ab0), .a2b1(din_23_ab1),
           .a2b0_1sc(din_23_ab0_1sc), .a2b1_1sc(din_23_ab1_1sc),
           .msk_a2b0(din_23_msk_ab0), .msk_a2b1(din_23_msk_ab1),
           .msk_a2b0_1sc(din_23_msk_ab0_1sc), .msk_a2b1_1sc(din_23_msk_ab1_1sc),
           
           .a3b0(din_25_ab0),
           .a3b0_1sc(din_25_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_20_calc (
           .clk(clk), .sign(din_signs_reg[20]), 
           .p(addr_7_20),
           .a0b0(din_20_ab0), .a0b1(din_20_ab1), .a0b2(din_20_ab2), .a0b3(din_20_ab3),
           .a0b0_1sc(din_20_ab0_1sc), .a0b1_1sc(din_20_ab1_1sc), .a0b2_1sc(din_20_ab2_1sc), .a0b3_1sc(din_20_ab3_1sc),
           .msk_a0b0(din_20_msk_ab0), .msk_a0b1(din_20_msk_ab1), .msk_a0b2(din_20_msk_ab2), .msk_a0b3(din_20_msk_ab3),
           .msk_a0b0_1sc(din_20_msk_ab0_1sc), .msk_a0b1_1sc(din_20_msk_ab1_1sc), .msk_a0b2_1sc(din_20_msk_ab2_1sc), .msk_a0b3_1sc(din_20_msk_ab3_1sc),

           .a1b0(din_22_ab0), .a1b1(din_22_ab1), .a1b2(din_22_ab2),
           .a1b0_1sc(din_22_ab0_1sc), .a1b1_1sc(din_22_ab1_1sc), .a1b2_1sc(din_22_ab2_1sc),
           .msk_a1b0(din_22_msk_ab0), .msk_a1b1(din_22_msk_ab1), .msk_a1b2(din_22_msk_ab2),
           .msk_a1b0_1sc(din_22_msk_ab0_1sc), .msk_a1b1_1sc(din_22_msk_ab1_1sc), .msk_a1b2_1sc(din_22_msk_ab2_1sc),

           .a2b0(din_24_ab0), .a2b1(din_24_ab1),
           .a2b0_1sc(din_24_ab0_1sc), .a2b1_1sc(din_24_ab1_1sc),
           .msk_a2b0(din_24_msk_ab0), .msk_a2b1(din_24_msk_ab1),
           .msk_a2b0_1sc(din_24_msk_ab0_1sc), .msk_a2b1_1sc(din_24_msk_ab1_1sc),
           
           .a3b0(din_26_ab0),
           .a3b0_1sc(din_26_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_21_calc (
           .clk(clk), .sign(din_signs_reg[21]), 
           .p(addr_7_21),
           .a0b0(din_21_ab0), .a0b1(din_21_ab1), .a0b2(din_21_ab2), .a0b3(din_21_ab3),
           .a0b0_1sc(din_21_ab0_1sc), .a0b1_1sc(din_21_ab1_1sc), .a0b2_1sc(din_21_ab2_1sc), .a0b3_1sc(din_21_ab3_1sc),
           .msk_a0b0(din_21_msk_ab0), .msk_a0b1(din_21_msk_ab1), .msk_a0b2(din_21_msk_ab2), .msk_a0b3(din_21_msk_ab3),
           .msk_a0b0_1sc(din_21_msk_ab0_1sc), .msk_a0b1_1sc(din_21_msk_ab1_1sc), .msk_a0b2_1sc(din_21_msk_ab2_1sc), .msk_a0b3_1sc(din_21_msk_ab3_1sc),

           .a1b0(din_23_ab0), .a1b1(din_23_ab1), .a1b2(din_23_ab2),
           .a1b0_1sc(din_23_ab0_1sc), .a1b1_1sc(din_23_ab1_1sc), .a1b2_1sc(din_23_ab2_1sc),
           .msk_a1b0(din_23_msk_ab0), .msk_a1b1(din_23_msk_ab1), .msk_a1b2(din_23_msk_ab2),
           .msk_a1b0_1sc(din_23_msk_ab0_1sc), .msk_a1b1_1sc(din_23_msk_ab1_1sc), .msk_a1b2_1sc(din_23_msk_ab2_1sc),

           .a2b0(din_25_ab0), .a2b1(din_25_ab1),
           .a2b0_1sc(din_25_ab0_1sc), .a2b1_1sc(din_25_ab1_1sc),
           .msk_a2b0(din_25_msk_ab0), .msk_a2b1(din_25_msk_ab1),
           .msk_a2b0_1sc(din_25_msk_ab0_1sc), .msk_a2b1_1sc(din_25_msk_ab1_1sc),
           
           .a3b0(din_27_ab0),
           .a3b0_1sc(din_27_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_22_calc (
           .clk(clk), .sign(din_signs_reg[22]), 
           .p(addr_7_22),
           .a0b0(din_22_ab0), .a0b1(din_22_ab1), .a0b2(din_22_ab2), .a0b3(din_22_ab3),
           .a0b0_1sc(din_22_ab0_1sc), .a0b1_1sc(din_22_ab1_1sc), .a0b2_1sc(din_22_ab2_1sc), .a0b3_1sc(din_22_ab3_1sc),
           .msk_a0b0(din_22_msk_ab0), .msk_a0b1(din_22_msk_ab1), .msk_a0b2(din_22_msk_ab2), .msk_a0b3(din_22_msk_ab3),
           .msk_a0b0_1sc(din_22_msk_ab0_1sc), .msk_a0b1_1sc(din_22_msk_ab1_1sc), .msk_a0b2_1sc(din_22_msk_ab2_1sc), .msk_a0b3_1sc(din_22_msk_ab3_1sc),

           .a1b0(din_24_ab0), .a1b1(din_24_ab1), .a1b2(din_24_ab2),
           .a1b0_1sc(din_24_ab0_1sc), .a1b1_1sc(din_24_ab1_1sc), .a1b2_1sc(din_24_ab2_1sc),
           .msk_a1b0(din_24_msk_ab0), .msk_a1b1(din_24_msk_ab1), .msk_a1b2(din_24_msk_ab2),
           .msk_a1b0_1sc(din_24_msk_ab0_1sc), .msk_a1b1_1sc(din_24_msk_ab1_1sc), .msk_a1b2_1sc(din_24_msk_ab2_1sc),

           .a2b0(din_26_ab0), .a2b1(din_26_ab1),
           .a2b0_1sc(din_26_ab0_1sc), .a2b1_1sc(din_26_ab1_1sc),
           .msk_a2b0(din_26_msk_ab0), .msk_a2b1(din_26_msk_ab1),
           .msk_a2b0_1sc(din_26_msk_ab0_1sc), .msk_a2b1_1sc(din_26_msk_ab1_1sc),
           
           .a3b0(din_28_ab0),
           .a3b0_1sc(din_28_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_23_calc (
           .clk(clk), .sign(din_signs_reg[23]), 
           .p(addr_7_23),
           .a0b0(din_23_ab0), .a0b1(din_23_ab1), .a0b2(din_23_ab2), .a0b3(din_23_ab3),
           .a0b0_1sc(din_23_ab0_1sc), .a0b1_1sc(din_23_ab1_1sc), .a0b2_1sc(din_23_ab2_1sc), .a0b3_1sc(din_23_ab3_1sc),
           .msk_a0b0(din_23_msk_ab0), .msk_a0b1(din_23_msk_ab1), .msk_a0b2(din_23_msk_ab2), .msk_a0b3(din_23_msk_ab3),
           .msk_a0b0_1sc(din_23_msk_ab0_1sc), .msk_a0b1_1sc(din_23_msk_ab1_1sc), .msk_a0b2_1sc(din_23_msk_ab2_1sc), .msk_a0b3_1sc(din_23_msk_ab3_1sc),

           .a1b0(din_25_ab0), .a1b1(din_25_ab1), .a1b2(din_25_ab2),
           .a1b0_1sc(din_25_ab0_1sc), .a1b1_1sc(din_25_ab1_1sc), .a1b2_1sc(din_25_ab2_1sc),
           .msk_a1b0(din_25_msk_ab0), .msk_a1b1(din_25_msk_ab1), .msk_a1b2(din_25_msk_ab2),
           .msk_a1b0_1sc(din_25_msk_ab0_1sc), .msk_a1b1_1sc(din_25_msk_ab1_1sc), .msk_a1b2_1sc(din_25_msk_ab2_1sc),

           .a2b0(din_27_ab0), .a2b1(din_27_ab1),
           .a2b0_1sc(din_27_ab0_1sc), .a2b1_1sc(din_27_ab1_1sc),
           .msk_a2b0(din_27_msk_ab0), .msk_a2b1(din_27_msk_ab1),
           .msk_a2b0_1sc(din_27_msk_ab0_1sc), .msk_a2b1_1sc(din_27_msk_ab1_1sc),
           
           .a3b0(din_29_ab0),
           .a3b0_1sc(din_29_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_24_calc (
           .clk(clk), .sign(din_signs_reg[24]), 
           .p(addr_7_24),
           .a0b0(din_24_ab0), .a0b1(din_24_ab1), .a0b2(din_24_ab2), .a0b3(din_24_ab3),
           .a0b0_1sc(din_24_ab0_1sc), .a0b1_1sc(din_24_ab1_1sc), .a0b2_1sc(din_24_ab2_1sc), .a0b3_1sc(din_24_ab3_1sc),
           .msk_a0b0(din_24_msk_ab0), .msk_a0b1(din_24_msk_ab1), .msk_a0b2(din_24_msk_ab2), .msk_a0b3(din_24_msk_ab3),
           .msk_a0b0_1sc(din_24_msk_ab0_1sc), .msk_a0b1_1sc(din_24_msk_ab1_1sc), .msk_a0b2_1sc(din_24_msk_ab2_1sc), .msk_a0b3_1sc(din_24_msk_ab3_1sc),

           .a1b0(din_26_ab0), .a1b1(din_26_ab1), .a1b2(din_26_ab2),
           .a1b0_1sc(din_26_ab0_1sc), .a1b1_1sc(din_26_ab1_1sc), .a1b2_1sc(din_26_ab2_1sc),
           .msk_a1b0(din_26_msk_ab0), .msk_a1b1(din_26_msk_ab1), .msk_a1b2(din_26_msk_ab2),
           .msk_a1b0_1sc(din_26_msk_ab0_1sc), .msk_a1b1_1sc(din_26_msk_ab1_1sc), .msk_a1b2_1sc(din_26_msk_ab2_1sc),

           .a2b0(din_28_ab0), .a2b1(din_28_ab1),
           .a2b0_1sc(din_28_ab0_1sc), .a2b1_1sc(din_28_ab1_1sc),
           .msk_a2b0(din_28_msk_ab0), .msk_a2b1(din_28_msk_ab1),
           .msk_a2b0_1sc(din_28_msk_ab0_1sc), .msk_a2b1_1sc(din_28_msk_ab1_1sc),
           
           .a3b0(din_30_ab0),
           .a3b0_1sc(din_30_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_25_calc (
           .clk(clk), .sign(din_signs_reg[25]), 
           .p(addr_7_25),
           .a0b0(din_25_ab0), .a0b1(din_25_ab1), .a0b2(din_25_ab2), .a0b3(din_25_ab3),
           .a0b0_1sc(din_25_ab0_1sc), .a0b1_1sc(din_25_ab1_1sc), .a0b2_1sc(din_25_ab2_1sc), .a0b3_1sc(din_25_ab3_1sc),
           .msk_a0b0(din_25_msk_ab0), .msk_a0b1(din_25_msk_ab1), .msk_a0b2(din_25_msk_ab2), .msk_a0b3(din_25_msk_ab3),
           .msk_a0b0_1sc(din_25_msk_ab0_1sc), .msk_a0b1_1sc(din_25_msk_ab1_1sc), .msk_a0b2_1sc(din_25_msk_ab2_1sc), .msk_a0b3_1sc(din_25_msk_ab3_1sc),

           .a1b0(din_27_ab0), .a1b1(din_27_ab1), .a1b2(din_27_ab2),
           .a1b0_1sc(din_27_ab0_1sc), .a1b1_1sc(din_27_ab1_1sc), .a1b2_1sc(din_27_ab2_1sc),
           .msk_a1b0(din_27_msk_ab0), .msk_a1b1(din_27_msk_ab1), .msk_a1b2(din_27_msk_ab2),
           .msk_a1b0_1sc(din_27_msk_ab0_1sc), .msk_a1b1_1sc(din_27_msk_ab1_1sc), .msk_a1b2_1sc(din_27_msk_ab2_1sc),

           .a2b0(din_29_ab0), .a2b1(din_29_ab1),
           .a2b0_1sc(din_29_ab0_1sc), .a2b1_1sc(din_29_ab1_1sc),
           .msk_a2b0(din_29_msk_ab0), .msk_a2b1(din_29_msk_ab1),
           .msk_a2b0_1sc(din_29_msk_ab0_1sc), .msk_a2b1_1sc(din_29_msk_ab1_1sc),
           
           .a3b0(din_31_ab0),
           .a3b0_1sc(din_31_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_26_calc (
           .clk(clk), .sign(din_signs_reg[26]), 
           .p(addr_7_26),
           .a0b0(din_26_ab0), .a0b1(din_26_ab1), .a0b2(din_26_ab2), .a0b3(din_26_ab3),
           .a0b0_1sc(din_26_ab0_1sc), .a0b1_1sc(din_26_ab1_1sc), .a0b2_1sc(din_26_ab2_1sc), .a0b3_1sc(din_26_ab3_1sc),
           .msk_a0b0(din_26_msk_ab0), .msk_a0b1(din_26_msk_ab1), .msk_a0b2(din_26_msk_ab2), .msk_a0b3(din_26_msk_ab3),
           .msk_a0b0_1sc(din_26_msk_ab0_1sc), .msk_a0b1_1sc(din_26_msk_ab1_1sc), .msk_a0b2_1sc(din_26_msk_ab2_1sc), .msk_a0b3_1sc(din_26_msk_ab3_1sc),

           .a1b0(din_28_ab0), .a1b1(din_28_ab1), .a1b2(din_28_ab2),
           .a1b0_1sc(din_28_ab0_1sc), .a1b1_1sc(din_28_ab1_1sc), .a1b2_1sc(din_28_ab2_1sc),
           .msk_a1b0(din_28_msk_ab0), .msk_a1b1(din_28_msk_ab1), .msk_a1b2(din_28_msk_ab2),
           .msk_a1b0_1sc(din_28_msk_ab0_1sc), .msk_a1b1_1sc(din_28_msk_ab1_1sc), .msk_a1b2_1sc(din_28_msk_ab2_1sc),

           .a2b0(din_30_ab0), .a2b1(din_30_ab1),
           .a2b0_1sc(din_30_ab0_1sc), .a2b1_1sc(din_30_ab1_1sc),
           .msk_a2b0(din_30_msk_ab0), .msk_a2b1(din_30_msk_ab1),
           .msk_a2b0_1sc(din_30_msk_ab0_1sc), .msk_a2b1_1sc(din_30_msk_ab1_1sc),
           
           .a3b0(din_32_ab0),
           .a3b0_1sc(din_32_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_27_calc (
           .clk(clk), .sign(din_signs_reg[27]), 
           .p(addr_7_27),
           .a0b0(din_27_ab0), .a0b1(din_27_ab1), .a0b2(din_27_ab2), .a0b3(din_27_ab3),
           .a0b0_1sc(din_27_ab0_1sc), .a0b1_1sc(din_27_ab1_1sc), .a0b2_1sc(din_27_ab2_1sc), .a0b3_1sc(din_27_ab3_1sc),
           .msk_a0b0(din_27_msk_ab0), .msk_a0b1(din_27_msk_ab1), .msk_a0b2(din_27_msk_ab2), .msk_a0b3(din_27_msk_ab3),
           .msk_a0b0_1sc(din_27_msk_ab0_1sc), .msk_a0b1_1sc(din_27_msk_ab1_1sc), .msk_a0b2_1sc(din_27_msk_ab2_1sc), .msk_a0b3_1sc(din_27_msk_ab3_1sc),

           .a1b0(din_29_ab0), .a1b1(din_29_ab1), .a1b2(din_29_ab2),
           .a1b0_1sc(din_29_ab0_1sc), .a1b1_1sc(din_29_ab1_1sc), .a1b2_1sc(din_29_ab2_1sc),
           .msk_a1b0(din_29_msk_ab0), .msk_a1b1(din_29_msk_ab1), .msk_a1b2(din_29_msk_ab2),
           .msk_a1b0_1sc(din_29_msk_ab0_1sc), .msk_a1b1_1sc(din_29_msk_ab1_1sc), .msk_a1b2_1sc(din_29_msk_ab2_1sc),

           .a2b0(din_31_ab0), .a2b1(din_31_ab1),
           .a2b0_1sc(din_31_ab0_1sc), .a2b1_1sc(din_31_ab1_1sc),
           .msk_a2b0(din_31_msk_ab0), .msk_a2b1(din_31_msk_ab1),
           .msk_a2b0_1sc(din_31_msk_ab0_1sc), .msk_a2b1_1sc(din_31_msk_ab1_1sc),
           
           .a3b0(din_33_ab0),
           .a3b0_1sc(din_33_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_28_calc (
           .clk(clk), .sign(din_signs_reg[28]), 
           .p(addr_7_28),
           .a0b0(din_28_ab0), .a0b1(din_28_ab1), .a0b2(din_28_ab2), .a0b3(din_28_ab3),
           .a0b0_1sc(din_28_ab0_1sc), .a0b1_1sc(din_28_ab1_1sc), .a0b2_1sc(din_28_ab2_1sc), .a0b3_1sc(din_28_ab3_1sc),
           .msk_a0b0(din_28_msk_ab0), .msk_a0b1(din_28_msk_ab1), .msk_a0b2(din_28_msk_ab2), .msk_a0b3(din_28_msk_ab3),
           .msk_a0b0_1sc(din_28_msk_ab0_1sc), .msk_a0b1_1sc(din_28_msk_ab1_1sc), .msk_a0b2_1sc(din_28_msk_ab2_1sc), .msk_a0b3_1sc(din_28_msk_ab3_1sc),

           .a1b0(din_30_ab0), .a1b1(din_30_ab1), .a1b2(din_30_ab2),
           .a1b0_1sc(din_30_ab0_1sc), .a1b1_1sc(din_30_ab1_1sc), .a1b2_1sc(din_30_ab2_1sc),
           .msk_a1b0(din_30_msk_ab0), .msk_a1b1(din_30_msk_ab1), .msk_a1b2(din_30_msk_ab2),
           .msk_a1b0_1sc(din_30_msk_ab0_1sc), .msk_a1b1_1sc(din_30_msk_ab1_1sc), .msk_a1b2_1sc(din_30_msk_ab2_1sc),

           .a2b0(din_32_ab0), .a2b1(din_32_ab1),
           .a2b0_1sc(din_32_ab0_1sc), .a2b1_1sc(din_32_ab1_1sc),
           .msk_a2b0(din_32_msk_ab0), .msk_a2b1(din_32_msk_ab1),
           .msk_a2b0_1sc(din_32_msk_ab0_1sc), .msk_a2b1_1sc(din_32_msk_ab1_1sc),
           
           .a3b0(din_34_ab0),
           .a3b0_1sc(din_34_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_29_calc (
           .clk(clk), .sign(din_signs_reg[29]), 
           .p(addr_7_29),
           .a0b0(din_29_ab0), .a0b1(din_29_ab1), .a0b2(din_29_ab2), .a0b3(din_29_ab3),
           .a0b0_1sc(din_29_ab0_1sc), .a0b1_1sc(din_29_ab1_1sc), .a0b2_1sc(din_29_ab2_1sc), .a0b3_1sc(din_29_ab3_1sc),
           .msk_a0b0(din_29_msk_ab0), .msk_a0b1(din_29_msk_ab1), .msk_a0b2(din_29_msk_ab2), .msk_a0b3(din_29_msk_ab3),
           .msk_a0b0_1sc(din_29_msk_ab0_1sc), .msk_a0b1_1sc(din_29_msk_ab1_1sc), .msk_a0b2_1sc(din_29_msk_ab2_1sc), .msk_a0b3_1sc(din_29_msk_ab3_1sc),

           .a1b0(din_31_ab0), .a1b1(din_31_ab1), .a1b2(din_31_ab2),
           .a1b0_1sc(din_31_ab0_1sc), .a1b1_1sc(din_31_ab1_1sc), .a1b2_1sc(din_31_ab2_1sc),
           .msk_a1b0(din_31_msk_ab0), .msk_a1b1(din_31_msk_ab1), .msk_a1b2(din_31_msk_ab2),
           .msk_a1b0_1sc(din_31_msk_ab0_1sc), .msk_a1b1_1sc(din_31_msk_ab1_1sc), .msk_a1b2_1sc(din_31_msk_ab2_1sc),

           .a2b0(din_33_ab0), .a2b1(din_33_ab1),
           .a2b0_1sc(din_33_ab0_1sc), .a2b1_1sc(din_33_ab1_1sc),
           .msk_a2b0(din_33_msk_ab0), .msk_a2b1(din_33_msk_ab1),
           .msk_a2b0_1sc(din_33_msk_ab0_1sc), .msk_a2b1_1sc(din_33_msk_ab1_1sc),
           
           .a3b0(din_35_ab0),
           .a3b0_1sc(din_35_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_30_calc (
           .clk(clk), .sign(din_signs_reg[30]), 
           .p(addr_7_30),
           .a0b0(din_30_ab0), .a0b1(din_30_ab1), .a0b2(din_30_ab2), .a0b3(din_30_ab3),
           .a0b0_1sc(din_30_ab0_1sc), .a0b1_1sc(din_30_ab1_1sc), .a0b2_1sc(din_30_ab2_1sc), .a0b3_1sc(din_30_ab3_1sc),
           .msk_a0b0(din_30_msk_ab0), .msk_a0b1(din_30_msk_ab1), .msk_a0b2(din_30_msk_ab2), .msk_a0b3(din_30_msk_ab3),
           .msk_a0b0_1sc(din_30_msk_ab0_1sc), .msk_a0b1_1sc(din_30_msk_ab1_1sc), .msk_a0b2_1sc(din_30_msk_ab2_1sc), .msk_a0b3_1sc(din_30_msk_ab3_1sc),

           .a1b0(din_32_ab0), .a1b1(din_32_ab1), .a1b2(din_32_ab2),
           .a1b0_1sc(din_32_ab0_1sc), .a1b1_1sc(din_32_ab1_1sc), .a1b2_1sc(din_32_ab2_1sc),
           .msk_a1b0(din_32_msk_ab0), .msk_a1b1(din_32_msk_ab1), .msk_a1b2(din_32_msk_ab2),
           .msk_a1b0_1sc(din_32_msk_ab0_1sc), .msk_a1b1_1sc(din_32_msk_ab1_1sc), .msk_a1b2_1sc(din_32_msk_ab2_1sc),

           .a2b0(din_34_ab0), .a2b1(din_34_ab1),
           .a2b0_1sc(din_34_ab0_1sc), .a2b1_1sc(din_34_ab1_1sc),
           .msk_a2b0(din_34_msk_ab0), .msk_a2b1(din_34_msk_ab1),
           .msk_a2b0_1sc(din_34_msk_ab0_1sc), .msk_a2b1_1sc(din_34_msk_ab1_1sc),
           
           .a3b0(din_36_ab0),
           .a3b0_1sc(din_36_ab0_1sc)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(8)
) addr_7_31_calc (
           .clk(clk), .sign(din_signs_reg[31]), 
           .p(addr_7_31),
           .a0b0(din_31_ab0), .a0b1(din_31_ab1), .a0b2(din_31_ab2), .a0b3(din_31_ab3),
           .a0b0_1sc(din_31_ab0_1sc), .a0b1_1sc(din_31_ab1_1sc), .a0b2_1sc(din_31_ab2_1sc), .a0b3_1sc(din_31_ab3_1sc),
           .msk_a0b0(din_31_msk_ab0), .msk_a0b1(din_31_msk_ab1), .msk_a0b2(din_31_msk_ab2), .msk_a0b3(din_31_msk_ab3),
           .msk_a0b0_1sc(din_31_msk_ab0_1sc), .msk_a0b1_1sc(din_31_msk_ab1_1sc), .msk_a0b2_1sc(din_31_msk_ab2_1sc), .msk_a0b3_1sc(din_31_msk_ab3_1sc),

           .a1b0(din_33_ab0), .a1b1(din_33_ab1), .a1b2(din_33_ab2),
           .a1b0_1sc(din_33_ab0_1sc), .a1b1_1sc(din_33_ab1_1sc), .a1b2_1sc(din_33_ab2_1sc),
           .msk_a1b0(din_33_msk_ab0), .msk_a1b1(din_33_msk_ab1), .msk_a1b2(din_33_msk_ab2),
           .msk_a1b0_1sc(din_33_msk_ab0_1sc), .msk_a1b1_1sc(din_33_msk_ab1_1sc), .msk_a1b2_1sc(din_33_msk_ab2_1sc),

           .a2b0(din_35_ab0), .a2b1(din_35_ab1),
           .a2b0_1sc(din_35_ab0_1sc), .a2b1_1sc(din_35_ab1_1sc),
           .msk_a2b0(din_35_msk_ab0), .msk_a2b1(din_35_msk_ab1),
           .msk_a2b0_1sc(din_35_msk_ab0_1sc), .msk_a2b1_1sc(din_35_msk_ab1_1sc),
           
           .a3b0(din_37_ab0),
           .a3b0_1sc(din_37_ab0_1sc)
);



hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_0 (
	.clk (clk),
	.addr0 (addr_0_0),
	.addr0_valid (addr_valid_0_0),
	.addr1 (addr_0_1),
	.addr1_valid (addr_valid_0_1),
	.dout0 (dout_0_0),
	.dout0_valid (dout_valid_0_0),
	.dout1 (dout_0_1),
	.dout1_valid (dout_valid_0_1)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_1 (
	.clk (clk),
	.addr0 (addr_0_2),
	.addr0_valid (addr_valid_0_2),
	.addr1 (addr_0_3),
	.addr1_valid (addr_valid_0_3),
	.dout0 (dout_0_2),
	.dout0_valid (dout_valid_0_2),
	.dout1 (dout_0_3),
	.dout1_valid (dout_valid_0_3)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_2 (
	.clk (clk),
	.addr0 (addr_0_4),
	.addr0_valid (addr_valid_0_4),
	.addr1 (addr_0_5),
	.addr1_valid (addr_valid_0_5),
	.dout0 (dout_0_4),
	.dout0_valid (dout_valid_0_4),
	.dout1 (dout_0_5),
	.dout1_valid (dout_valid_0_5)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_3 (
	.clk (clk),
	.addr0 (addr_0_6),
	.addr0_valid (addr_valid_0_6),
	.addr1 (addr_0_7),
	.addr1_valid (addr_valid_0_7),
	.dout0 (dout_0_6),
	.dout0_valid (dout_valid_0_6),
	.dout1 (dout_0_7),
	.dout1_valid (dout_valid_0_7)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_4 (
	.clk (clk),
	.addr0 (addr_0_8),
	.addr0_valid (addr_valid_0_8),
	.addr1 (addr_0_9),
	.addr1_valid (addr_valid_0_9),
	.dout0 (dout_0_8),
	.dout0_valid (dout_valid_0_8),
	.dout1 (dout_0_9),
	.dout1_valid (dout_valid_0_9)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_5 (
	.clk (clk),
	.addr0 (addr_0_10),
	.addr0_valid (addr_valid_0_10),
	.addr1 (addr_0_11),
	.addr1_valid (addr_valid_0_11),
	.dout0 (dout_0_10),
	.dout0_valid (dout_valid_0_10),
	.dout1 (dout_0_11),
	.dout1_valid (dout_valid_0_11)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_6 (
	.clk (clk),
	.addr0 (addr_0_12),
	.addr0_valid (addr_valid_0_12),
	.addr1 (addr_0_13),
	.addr1_valid (addr_valid_0_13),
	.dout0 (dout_0_12),
	.dout0_valid (dout_valid_0_12),
	.dout1 (dout_0_13),
	.dout1_valid (dout_valid_0_13)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_7 (
	.clk (clk),
	.addr0 (addr_0_14),
	.addr0_valid (addr_valid_0_14),
	.addr1 (addr_0_15),
	.addr1_valid (addr_valid_0_15),
	.dout0 (dout_0_14),
	.dout0_valid (dout_valid_0_14),
	.dout1 (dout_0_15),
	.dout1_valid (dout_valid_0_15)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_8 (
	.clk (clk),
	.addr0 (addr_0_16),
	.addr0_valid (addr_valid_0_16),
	.addr1 (addr_0_17),
	.addr1_valid (addr_valid_0_17),
	.dout0 (dout_0_16),
	.dout0_valid (dout_valid_0_16),
	.dout1 (dout_0_17),
	.dout1_valid (dout_valid_0_17)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_9 (
	.clk (clk),
	.addr0 (addr_0_18),
	.addr0_valid (addr_valid_0_18),
	.addr1 (addr_0_19),
	.addr1_valid (addr_valid_0_19),
	.dout0 (dout_0_18),
	.dout0_valid (dout_valid_0_18),
	.dout1 (dout_0_19),
	.dout1_valid (dout_valid_0_19)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_10 (
	.clk (clk),
	.addr0 (addr_0_20),
	.addr0_valid (addr_valid_0_20),
	.addr1 (addr_0_21),
	.addr1_valid (addr_valid_0_21),
	.dout0 (dout_0_20),
	.dout0_valid (dout_valid_0_20),
	.dout1 (dout_0_21),
	.dout1_valid (dout_valid_0_21)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_11 (
	.clk (clk),
	.addr0 (addr_0_22),
	.addr0_valid (addr_valid_0_22),
	.addr1 (addr_0_23),
	.addr1_valid (addr_valid_0_23),
	.dout0 (dout_0_22),
	.dout0_valid (dout_valid_0_22),
	.dout1 (dout_0_23),
	.dout1_valid (dout_valid_0_23)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_12 (
	.clk (clk),
	.addr0 (addr_0_24),
	.addr0_valid (addr_valid_0_24),
	.addr1 (addr_0_25),
	.addr1_valid (addr_valid_0_25),
	.dout0 (dout_0_24),
	.dout0_valid (dout_valid_0_24),
	.dout1 (dout_0_25),
	.dout1_valid (dout_valid_0_25)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_13 (
	.clk (clk),
	.addr0 (addr_0_26),
	.addr0_valid (addr_valid_0_26),
	.addr1 (addr_0_27),
	.addr1_valid (addr_valid_0_27),
	.dout0 (dout_0_26),
	.dout0_valid (dout_valid_0_26),
	.dout1 (dout_0_27),
	.dout1_valid (dout_valid_0_27)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_14 (
	.clk (clk),
	.addr0 (addr_0_28),
	.addr0_valid (addr_valid_0_28),
	.addr1 (addr_0_29),
	.addr1_valid (addr_valid_0_29),
	.dout0 (dout_0_28),
	.dout0_valid (dout_valid_0_28),
	.dout1 (dout_0_29),
	.dout1_valid (dout_valid_0_29)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap0.mif")
)
hashtable_0_15 (
	.clk (clk),
	.addr0 (addr_0_30),
	.addr0_valid (addr_valid_0_30),
	.addr1 (addr_0_31),
	.addr1_valid (addr_valid_0_31),
	.dout0 (dout_0_30),
	.dout0_valid (dout_valid_0_30),
	.dout1 (dout_0_31),
	.dout1_valid (dout_valid_0_31)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_0 (
	.clk (clk),
	.addr0 (addr_1_0),
	.addr0_valid (addr_valid_1_0),
	.addr1 (addr_1_1),
	.addr1_valid (addr_valid_1_1),
	.dout0 (dout_1_0),
	.dout0_valid (dout_valid_1_0),
	.dout1 (dout_1_1),
	.dout1_valid (dout_valid_1_1)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_1 (
	.clk (clk),
	.addr0 (addr_1_2),
	.addr0_valid (addr_valid_1_2),
	.addr1 (addr_1_3),
	.addr1_valid (addr_valid_1_3),
	.dout0 (dout_1_2),
	.dout0_valid (dout_valid_1_2),
	.dout1 (dout_1_3),
	.dout1_valid (dout_valid_1_3)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_2 (
	.clk (clk),
	.addr0 (addr_1_4),
	.addr0_valid (addr_valid_1_4),
	.addr1 (addr_1_5),
	.addr1_valid (addr_valid_1_5),
	.dout0 (dout_1_4),
	.dout0_valid (dout_valid_1_4),
	.dout1 (dout_1_5),
	.dout1_valid (dout_valid_1_5)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_3 (
	.clk (clk),
	.addr0 (addr_1_6),
	.addr0_valid (addr_valid_1_6),
	.addr1 (addr_1_7),
	.addr1_valid (addr_valid_1_7),
	.dout0 (dout_1_6),
	.dout0_valid (dout_valid_1_6),
	.dout1 (dout_1_7),
	.dout1_valid (dout_valid_1_7)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_4 (
	.clk (clk),
	.addr0 (addr_1_8),
	.addr0_valid (addr_valid_1_8),
	.addr1 (addr_1_9),
	.addr1_valid (addr_valid_1_9),
	.dout0 (dout_1_8),
	.dout0_valid (dout_valid_1_8),
	.dout1 (dout_1_9),
	.dout1_valid (dout_valid_1_9)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_5 (
	.clk (clk),
	.addr0 (addr_1_10),
	.addr0_valid (addr_valid_1_10),
	.addr1 (addr_1_11),
	.addr1_valid (addr_valid_1_11),
	.dout0 (dout_1_10),
	.dout0_valid (dout_valid_1_10),
	.dout1 (dout_1_11),
	.dout1_valid (dout_valid_1_11)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_6 (
	.clk (clk),
	.addr0 (addr_1_12),
	.addr0_valid (addr_valid_1_12),
	.addr1 (addr_1_13),
	.addr1_valid (addr_valid_1_13),
	.dout0 (dout_1_12),
	.dout0_valid (dout_valid_1_12),
	.dout1 (dout_1_13),
	.dout1_valid (dout_valid_1_13)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_7 (
	.clk (clk),
	.addr0 (addr_1_14),
	.addr0_valid (addr_valid_1_14),
	.addr1 (addr_1_15),
	.addr1_valid (addr_valid_1_15),
	.dout0 (dout_1_14),
	.dout0_valid (dout_valid_1_14),
	.dout1 (dout_1_15),
	.dout1_valid (dout_valid_1_15)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_8 (
	.clk (clk),
	.addr0 (addr_1_16),
	.addr0_valid (addr_valid_1_16),
	.addr1 (addr_1_17),
	.addr1_valid (addr_valid_1_17),
	.dout0 (dout_1_16),
	.dout0_valid (dout_valid_1_16),
	.dout1 (dout_1_17),
	.dout1_valid (dout_valid_1_17)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_9 (
	.clk (clk),
	.addr0 (addr_1_18),
	.addr0_valid (addr_valid_1_18),
	.addr1 (addr_1_19),
	.addr1_valid (addr_valid_1_19),
	.dout0 (dout_1_18),
	.dout0_valid (dout_valid_1_18),
	.dout1 (dout_1_19),
	.dout1_valid (dout_valid_1_19)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_10 (
	.clk (clk),
	.addr0 (addr_1_20),
	.addr0_valid (addr_valid_1_20),
	.addr1 (addr_1_21),
	.addr1_valid (addr_valid_1_21),
	.dout0 (dout_1_20),
	.dout0_valid (dout_valid_1_20),
	.dout1 (dout_1_21),
	.dout1_valid (dout_valid_1_21)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_11 (
	.clk (clk),
	.addr0 (addr_1_22),
	.addr0_valid (addr_valid_1_22),
	.addr1 (addr_1_23),
	.addr1_valid (addr_valid_1_23),
	.dout0 (dout_1_22),
	.dout0_valid (dout_valid_1_22),
	.dout1 (dout_1_23),
	.dout1_valid (dout_valid_1_23)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_12 (
	.clk (clk),
	.addr0 (addr_1_24),
	.addr0_valid (addr_valid_1_24),
	.addr1 (addr_1_25),
	.addr1_valid (addr_valid_1_25),
	.dout0 (dout_1_24),
	.dout0_valid (dout_valid_1_24),
	.dout1 (dout_1_25),
	.dout1_valid (dout_valid_1_25)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_13 (
	.clk (clk),
	.addr0 (addr_1_26),
	.addr0_valid (addr_valid_1_26),
	.addr1 (addr_1_27),
	.addr1_valid (addr_valid_1_27),
	.dout0 (dout_1_26),
	.dout0_valid (dout_valid_1_26),
	.dout1 (dout_1_27),
	.dout1_valid (dout_valid_1_27)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_14 (
	.clk (clk),
	.addr0 (addr_1_28),
	.addr0_valid (addr_valid_1_28),
	.addr1 (addr_1_29),
	.addr1_valid (addr_valid_1_29),
	.dout0 (dout_1_28),
	.dout0_valid (dout_valid_1_28),
	.dout1 (dout_1_29),
	.dout1_valid (dout_valid_1_29)
);

hashtable #(
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./memory_init/bitmap1.mif")
)
hashtable_1_15 (
	.clk (clk),
	.addr0 (addr_1_30),
	.addr0_valid (addr_valid_1_30),
	.addr1 (addr_1_31),
	.addr1_valid (addr_valid_1_31),
	.dout0 (dout_1_30),
	.dout0_valid (dout_valid_1_30),
	.dout1 (dout_1_31),
	.dout1_valid (dout_valid_1_31)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_0 (
	.clk (clk),
	.addr0 (addr_2_0),
	.addr0_valid (addr_valid_2_0),
	.addr1 (addr_2_1),
	.addr1_valid (addr_valid_2_1),
	.dout0 (dout_2_0),
	.dout0_valid (dout_valid_2_0),
	.dout1 (dout_2_1),
	.dout1_valid (dout_valid_2_1)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_1 (
	.clk (clk),
	.addr0 (addr_2_2),
	.addr0_valid (addr_valid_2_2),
	.addr1 (addr_2_3),
	.addr1_valid (addr_valid_2_3),
	.dout0 (dout_2_2),
	.dout0_valid (dout_valid_2_2),
	.dout1 (dout_2_3),
	.dout1_valid (dout_valid_2_3)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_2 (
	.clk (clk),
	.addr0 (addr_2_4),
	.addr0_valid (addr_valid_2_4),
	.addr1 (addr_2_5),
	.addr1_valid (addr_valid_2_5),
	.dout0 (dout_2_4),
	.dout0_valid (dout_valid_2_4),
	.dout1 (dout_2_5),
	.dout1_valid (dout_valid_2_5)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_3 (
	.clk (clk),
	.addr0 (addr_2_6),
	.addr0_valid (addr_valid_2_6),
	.addr1 (addr_2_7),
	.addr1_valid (addr_valid_2_7),
	.dout0 (dout_2_6),
	.dout0_valid (dout_valid_2_6),
	.dout1 (dout_2_7),
	.dout1_valid (dout_valid_2_7)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_4 (
	.clk (clk),
	.addr0 (addr_2_8),
	.addr0_valid (addr_valid_2_8),
	.addr1 (addr_2_9),
	.addr1_valid (addr_valid_2_9),
	.dout0 (dout_2_8),
	.dout0_valid (dout_valid_2_8),
	.dout1 (dout_2_9),
	.dout1_valid (dout_valid_2_9)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_5 (
	.clk (clk),
	.addr0 (addr_2_10),
	.addr0_valid (addr_valid_2_10),
	.addr1 (addr_2_11),
	.addr1_valid (addr_valid_2_11),
	.dout0 (dout_2_10),
	.dout0_valid (dout_valid_2_10),
	.dout1 (dout_2_11),
	.dout1_valid (dout_valid_2_11)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_6 (
	.clk (clk),
	.addr0 (addr_2_12),
	.addr0_valid (addr_valid_2_12),
	.addr1 (addr_2_13),
	.addr1_valid (addr_valid_2_13),
	.dout0 (dout_2_12),
	.dout0_valid (dout_valid_2_12),
	.dout1 (dout_2_13),
	.dout1_valid (dout_valid_2_13)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_7 (
	.clk (clk),
	.addr0 (addr_2_14),
	.addr0_valid (addr_valid_2_14),
	.addr1 (addr_2_15),
	.addr1_valid (addr_valid_2_15),
	.dout0 (dout_2_14),
	.dout0_valid (dout_valid_2_14),
	.dout1 (dout_2_15),
	.dout1_valid (dout_valid_2_15)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_8 (
	.clk (clk),
	.addr0 (addr_2_16),
	.addr0_valid (addr_valid_2_16),
	.addr1 (addr_2_17),
	.addr1_valid (addr_valid_2_17),
	.dout0 (dout_2_16),
	.dout0_valid (dout_valid_2_16),
	.dout1 (dout_2_17),
	.dout1_valid (dout_valid_2_17)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_9 (
	.clk (clk),
	.addr0 (addr_2_18),
	.addr0_valid (addr_valid_2_18),
	.addr1 (addr_2_19),
	.addr1_valid (addr_valid_2_19),
	.dout0 (dout_2_18),
	.dout0_valid (dout_valid_2_18),
	.dout1 (dout_2_19),
	.dout1_valid (dout_valid_2_19)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_10 (
	.clk (clk),
	.addr0 (addr_2_20),
	.addr0_valid (addr_valid_2_20),
	.addr1 (addr_2_21),
	.addr1_valid (addr_valid_2_21),
	.dout0 (dout_2_20),
	.dout0_valid (dout_valid_2_20),
	.dout1 (dout_2_21),
	.dout1_valid (dout_valid_2_21)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_11 (
	.clk (clk),
	.addr0 (addr_2_22),
	.addr0_valid (addr_valid_2_22),
	.addr1 (addr_2_23),
	.addr1_valid (addr_valid_2_23),
	.dout0 (dout_2_22),
	.dout0_valid (dout_valid_2_22),
	.dout1 (dout_2_23),
	.dout1_valid (dout_valid_2_23)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_12 (
	.clk (clk),
	.addr0 (addr_2_24),
	.addr0_valid (addr_valid_2_24),
	.addr1 (addr_2_25),
	.addr1_valid (addr_valid_2_25),
	.dout0 (dout_2_24),
	.dout0_valid (dout_valid_2_24),
	.dout1 (dout_2_25),
	.dout1_valid (dout_valid_2_25)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_13 (
	.clk (clk),
	.addr0 (addr_2_26),
	.addr0_valid (addr_valid_2_26),
	.addr1 (addr_2_27),
	.addr1_valid (addr_valid_2_27),
	.dout0 (dout_2_26),
	.dout0_valid (dout_valid_2_26),
	.dout1 (dout_2_27),
	.dout1_valid (dout_valid_2_27)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_14 (
	.clk (clk),
	.addr0 (addr_2_28),
	.addr0_valid (addr_valid_2_28),
	.addr1 (addr_2_29),
	.addr1_valid (addr_valid_2_29),
	.dout0 (dout_2_28),
	.dout0_valid (dout_valid_2_28),
	.dout1 (dout_2_29),
	.dout1_valid (dout_valid_2_29)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap2.mif")
)
hashtable_2_15 (
	.clk (clk),
	.addr0 (addr_2_30),
	.addr0_valid (addr_valid_2_30),
	.addr1 (addr_2_31),
	.addr1_valid (addr_valid_2_31),
	.dout0 (dout_2_30),
	.dout0_valid (dout_valid_2_30),
	.dout1 (dout_2_31),
	.dout1_valid (dout_valid_2_31)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_0 (
	.clk (clk),
	.addr0 (addr_3_0),
	.addr0_valid (addr_valid_3_0),
	.addr1 (addr_3_1),
	.addr1_valid (addr_valid_3_1),
	.dout0 (dout_3_0),
	.dout0_valid (dout_valid_3_0),
	.dout1 (dout_3_1),
	.dout1_valid (dout_valid_3_1)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_1 (
	.clk (clk),
	.addr0 (addr_3_2),
	.addr0_valid (addr_valid_3_2),
	.addr1 (addr_3_3),
	.addr1_valid (addr_valid_3_3),
	.dout0 (dout_3_2),
	.dout0_valid (dout_valid_3_2),
	.dout1 (dout_3_3),
	.dout1_valid (dout_valid_3_3)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_2 (
	.clk (clk),
	.addr0 (addr_3_4),
	.addr0_valid (addr_valid_3_4),
	.addr1 (addr_3_5),
	.addr1_valid (addr_valid_3_5),
	.dout0 (dout_3_4),
	.dout0_valid (dout_valid_3_4),
	.dout1 (dout_3_5),
	.dout1_valid (dout_valid_3_5)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_3 (
	.clk (clk),
	.addr0 (addr_3_6),
	.addr0_valid (addr_valid_3_6),
	.addr1 (addr_3_7),
	.addr1_valid (addr_valid_3_7),
	.dout0 (dout_3_6),
	.dout0_valid (dout_valid_3_6),
	.dout1 (dout_3_7),
	.dout1_valid (dout_valid_3_7)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_4 (
	.clk (clk),
	.addr0 (addr_3_8),
	.addr0_valid (addr_valid_3_8),
	.addr1 (addr_3_9),
	.addr1_valid (addr_valid_3_9),
	.dout0 (dout_3_8),
	.dout0_valid (dout_valid_3_8),
	.dout1 (dout_3_9),
	.dout1_valid (dout_valid_3_9)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_5 (
	.clk (clk),
	.addr0 (addr_3_10),
	.addr0_valid (addr_valid_3_10),
	.addr1 (addr_3_11),
	.addr1_valid (addr_valid_3_11),
	.dout0 (dout_3_10),
	.dout0_valid (dout_valid_3_10),
	.dout1 (dout_3_11),
	.dout1_valid (dout_valid_3_11)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_6 (
	.clk (clk),
	.addr0 (addr_3_12),
	.addr0_valid (addr_valid_3_12),
	.addr1 (addr_3_13),
	.addr1_valid (addr_valid_3_13),
	.dout0 (dout_3_12),
	.dout0_valid (dout_valid_3_12),
	.dout1 (dout_3_13),
	.dout1_valid (dout_valid_3_13)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_7 (
	.clk (clk),
	.addr0 (addr_3_14),
	.addr0_valid (addr_valid_3_14),
	.addr1 (addr_3_15),
	.addr1_valid (addr_valid_3_15),
	.dout0 (dout_3_14),
	.dout0_valid (dout_valid_3_14),
	.dout1 (dout_3_15),
	.dout1_valid (dout_valid_3_15)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_8 (
	.clk (clk),
	.addr0 (addr_3_16),
	.addr0_valid (addr_valid_3_16),
	.addr1 (addr_3_17),
	.addr1_valid (addr_valid_3_17),
	.dout0 (dout_3_16),
	.dout0_valid (dout_valid_3_16),
	.dout1 (dout_3_17),
	.dout1_valid (dout_valid_3_17)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_9 (
	.clk (clk),
	.addr0 (addr_3_18),
	.addr0_valid (addr_valid_3_18),
	.addr1 (addr_3_19),
	.addr1_valid (addr_valid_3_19),
	.dout0 (dout_3_18),
	.dout0_valid (dout_valid_3_18),
	.dout1 (dout_3_19),
	.dout1_valid (dout_valid_3_19)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_10 (
	.clk (clk),
	.addr0 (addr_3_20),
	.addr0_valid (addr_valid_3_20),
	.addr1 (addr_3_21),
	.addr1_valid (addr_valid_3_21),
	.dout0 (dout_3_20),
	.dout0_valid (dout_valid_3_20),
	.dout1 (dout_3_21),
	.dout1_valid (dout_valid_3_21)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_11 (
	.clk (clk),
	.addr0 (addr_3_22),
	.addr0_valid (addr_valid_3_22),
	.addr1 (addr_3_23),
	.addr1_valid (addr_valid_3_23),
	.dout0 (dout_3_22),
	.dout0_valid (dout_valid_3_22),
	.dout1 (dout_3_23),
	.dout1_valid (dout_valid_3_23)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_12 (
	.clk (clk),
	.addr0 (addr_3_24),
	.addr0_valid (addr_valid_3_24),
	.addr1 (addr_3_25),
	.addr1_valid (addr_valid_3_25),
	.dout0 (dout_3_24),
	.dout0_valid (dout_valid_3_24),
	.dout1 (dout_3_25),
	.dout1_valid (dout_valid_3_25)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_13 (
	.clk (clk),
	.addr0 (addr_3_26),
	.addr0_valid (addr_valid_3_26),
	.addr1 (addr_3_27),
	.addr1_valid (addr_valid_3_27),
	.dout0 (dout_3_26),
	.dout0_valid (dout_valid_3_26),
	.dout1 (dout_3_27),
	.dout1_valid (dout_valid_3_27)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_14 (
	.clk (clk),
	.addr0 (addr_3_28),
	.addr0_valid (addr_valid_3_28),
	.addr1 (addr_3_29),
	.addr1_valid (addr_valid_3_29),
	.dout0 (dout_3_28),
	.dout0_valid (dout_valid_3_28),
	.dout1 (dout_3_29),
	.dout1_valid (dout_valid_3_29)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap3.mif")
)
hashtable_3_15 (
	.clk (clk),
	.addr0 (addr_3_30),
	.addr0_valid (addr_valid_3_30),
	.addr1 (addr_3_31),
	.addr1_valid (addr_valid_3_31),
	.dout0 (dout_3_30),
	.dout0_valid (dout_valid_3_30),
	.dout1 (dout_3_31),
	.dout1_valid (dout_valid_3_31)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_0 (
	.clk (clk),
	.addr0 (addr_4_0),
	.addr0_valid (addr_valid_4_0),
	.addr1 (addr_4_1),
	.addr1_valid (addr_valid_4_1),
	.dout0 (dout_4_0),
	.dout0_valid (dout_valid_4_0),
	.dout1 (dout_4_1),
	.dout1_valid (dout_valid_4_1)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_1 (
	.clk (clk),
	.addr0 (addr_4_2),
	.addr0_valid (addr_valid_4_2),
	.addr1 (addr_4_3),
	.addr1_valid (addr_valid_4_3),
	.dout0 (dout_4_2),
	.dout0_valid (dout_valid_4_2),
	.dout1 (dout_4_3),
	.dout1_valid (dout_valid_4_3)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_2 (
	.clk (clk),
	.addr0 (addr_4_4),
	.addr0_valid (addr_valid_4_4),
	.addr1 (addr_4_5),
	.addr1_valid (addr_valid_4_5),
	.dout0 (dout_4_4),
	.dout0_valid (dout_valid_4_4),
	.dout1 (dout_4_5),
	.dout1_valid (dout_valid_4_5)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_3 (
	.clk (clk),
	.addr0 (addr_4_6),
	.addr0_valid (addr_valid_4_6),
	.addr1 (addr_4_7),
	.addr1_valid (addr_valid_4_7),
	.dout0 (dout_4_6),
	.dout0_valid (dout_valid_4_6),
	.dout1 (dout_4_7),
	.dout1_valid (dout_valid_4_7)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_4 (
	.clk (clk),
	.addr0 (addr_4_8),
	.addr0_valid (addr_valid_4_8),
	.addr1 (addr_4_9),
	.addr1_valid (addr_valid_4_9),
	.dout0 (dout_4_8),
	.dout0_valid (dout_valid_4_8),
	.dout1 (dout_4_9),
	.dout1_valid (dout_valid_4_9)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_5 (
	.clk (clk),
	.addr0 (addr_4_10),
	.addr0_valid (addr_valid_4_10),
	.addr1 (addr_4_11),
	.addr1_valid (addr_valid_4_11),
	.dout0 (dout_4_10),
	.dout0_valid (dout_valid_4_10),
	.dout1 (dout_4_11),
	.dout1_valid (dout_valid_4_11)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_6 (
	.clk (clk),
	.addr0 (addr_4_12),
	.addr0_valid (addr_valid_4_12),
	.addr1 (addr_4_13),
	.addr1_valid (addr_valid_4_13),
	.dout0 (dout_4_12),
	.dout0_valid (dout_valid_4_12),
	.dout1 (dout_4_13),
	.dout1_valid (dout_valid_4_13)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_7 (
	.clk (clk),
	.addr0 (addr_4_14),
	.addr0_valid (addr_valid_4_14),
	.addr1 (addr_4_15),
	.addr1_valid (addr_valid_4_15),
	.dout0 (dout_4_14),
	.dout0_valid (dout_valid_4_14),
	.dout1 (dout_4_15),
	.dout1_valid (dout_valid_4_15)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_8 (
	.clk (clk),
	.addr0 (addr_4_16),
	.addr0_valid (addr_valid_4_16),
	.addr1 (addr_4_17),
	.addr1_valid (addr_valid_4_17),
	.dout0 (dout_4_16),
	.dout0_valid (dout_valid_4_16),
	.dout1 (dout_4_17),
	.dout1_valid (dout_valid_4_17)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_9 (
	.clk (clk),
	.addr0 (addr_4_18),
	.addr0_valid (addr_valid_4_18),
	.addr1 (addr_4_19),
	.addr1_valid (addr_valid_4_19),
	.dout0 (dout_4_18),
	.dout0_valid (dout_valid_4_18),
	.dout1 (dout_4_19),
	.dout1_valid (dout_valid_4_19)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_10 (
	.clk (clk),
	.addr0 (addr_4_20),
	.addr0_valid (addr_valid_4_20),
	.addr1 (addr_4_21),
	.addr1_valid (addr_valid_4_21),
	.dout0 (dout_4_20),
	.dout0_valid (dout_valid_4_20),
	.dout1 (dout_4_21),
	.dout1_valid (dout_valid_4_21)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_11 (
	.clk (clk),
	.addr0 (addr_4_22),
	.addr0_valid (addr_valid_4_22),
	.addr1 (addr_4_23),
	.addr1_valid (addr_valid_4_23),
	.dout0 (dout_4_22),
	.dout0_valid (dout_valid_4_22),
	.dout1 (dout_4_23),
	.dout1_valid (dout_valid_4_23)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_12 (
	.clk (clk),
	.addr0 (addr_4_24),
	.addr0_valid (addr_valid_4_24),
	.addr1 (addr_4_25),
	.addr1_valid (addr_valid_4_25),
	.dout0 (dout_4_24),
	.dout0_valid (dout_valid_4_24),
	.dout1 (dout_4_25),
	.dout1_valid (dout_valid_4_25)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_13 (
	.clk (clk),
	.addr0 (addr_4_26),
	.addr0_valid (addr_valid_4_26),
	.addr1 (addr_4_27),
	.addr1_valid (addr_valid_4_27),
	.dout0 (dout_4_26),
	.dout0_valid (dout_valid_4_26),
	.dout1 (dout_4_27),
	.dout1_valid (dout_valid_4_27)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_14 (
	.clk (clk),
	.addr0 (addr_4_28),
	.addr0_valid (addr_valid_4_28),
	.addr1 (addr_4_29),
	.addr1_valid (addr_valid_4_29),
	.dout0 (dout_4_28),
	.dout0_valid (dout_valid_4_28),
	.dout1 (dout_4_29),
	.dout1_valid (dout_valid_4_29)
);

hashtable #(
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./memory_init/bitmap4.mif")
)
hashtable_4_15 (
	.clk (clk),
	.addr0 (addr_4_30),
	.addr0_valid (addr_valid_4_30),
	.addr1 (addr_4_31),
	.addr1_valid (addr_valid_4_31),
	.dout0 (dout_4_30),
	.dout0_valid (dout_valid_4_30),
	.dout1 (dout_4_31),
	.dout1_valid (dout_valid_4_31)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_0 (
	.clk (clk),
	.addr0 (addr_5_0),
	.addr0_valid (addr_valid_5_0),
	.addr1 (addr_5_1),
	.addr1_valid (addr_valid_5_1),
	.dout0 (dout_5_0),
	.dout0_valid (dout_valid_5_0),
	.dout1 (dout_5_1),
	.dout1_valid (dout_valid_5_1)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_1 (
	.clk (clk),
	.addr0 (addr_5_2),
	.addr0_valid (addr_valid_5_2),
	.addr1 (addr_5_3),
	.addr1_valid (addr_valid_5_3),
	.dout0 (dout_5_2),
	.dout0_valid (dout_valid_5_2),
	.dout1 (dout_5_3),
	.dout1_valid (dout_valid_5_3)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_2 (
	.clk (clk),
	.addr0 (addr_5_4),
	.addr0_valid (addr_valid_5_4),
	.addr1 (addr_5_5),
	.addr1_valid (addr_valid_5_5),
	.dout0 (dout_5_4),
	.dout0_valid (dout_valid_5_4),
	.dout1 (dout_5_5),
	.dout1_valid (dout_valid_5_5)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_3 (
	.clk (clk),
	.addr0 (addr_5_6),
	.addr0_valid (addr_valid_5_6),
	.addr1 (addr_5_7),
	.addr1_valid (addr_valid_5_7),
	.dout0 (dout_5_6),
	.dout0_valid (dout_valid_5_6),
	.dout1 (dout_5_7),
	.dout1_valid (dout_valid_5_7)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_4 (
	.clk (clk),
	.addr0 (addr_5_8),
	.addr0_valid (addr_valid_5_8),
	.addr1 (addr_5_9),
	.addr1_valid (addr_valid_5_9),
	.dout0 (dout_5_8),
	.dout0_valid (dout_valid_5_8),
	.dout1 (dout_5_9),
	.dout1_valid (dout_valid_5_9)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_5 (
	.clk (clk),
	.addr0 (addr_5_10),
	.addr0_valid (addr_valid_5_10),
	.addr1 (addr_5_11),
	.addr1_valid (addr_valid_5_11),
	.dout0 (dout_5_10),
	.dout0_valid (dout_valid_5_10),
	.dout1 (dout_5_11),
	.dout1_valid (dout_valid_5_11)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_6 (
	.clk (clk),
	.addr0 (addr_5_12),
	.addr0_valid (addr_valid_5_12),
	.addr1 (addr_5_13),
	.addr1_valid (addr_valid_5_13),
	.dout0 (dout_5_12),
	.dout0_valid (dout_valid_5_12),
	.dout1 (dout_5_13),
	.dout1_valid (dout_valid_5_13)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_7 (
	.clk (clk),
	.addr0 (addr_5_14),
	.addr0_valid (addr_valid_5_14),
	.addr1 (addr_5_15),
	.addr1_valid (addr_valid_5_15),
	.dout0 (dout_5_14),
	.dout0_valid (dout_valid_5_14),
	.dout1 (dout_5_15),
	.dout1_valid (dout_valid_5_15)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_8 (
	.clk (clk),
	.addr0 (addr_5_16),
	.addr0_valid (addr_valid_5_16),
	.addr1 (addr_5_17),
	.addr1_valid (addr_valid_5_17),
	.dout0 (dout_5_16),
	.dout0_valid (dout_valid_5_16),
	.dout1 (dout_5_17),
	.dout1_valid (dout_valid_5_17)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_9 (
	.clk (clk),
	.addr0 (addr_5_18),
	.addr0_valid (addr_valid_5_18),
	.addr1 (addr_5_19),
	.addr1_valid (addr_valid_5_19),
	.dout0 (dout_5_18),
	.dout0_valid (dout_valid_5_18),
	.dout1 (dout_5_19),
	.dout1_valid (dout_valid_5_19)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_10 (
	.clk (clk),
	.addr0 (addr_5_20),
	.addr0_valid (addr_valid_5_20),
	.addr1 (addr_5_21),
	.addr1_valid (addr_valid_5_21),
	.dout0 (dout_5_20),
	.dout0_valid (dout_valid_5_20),
	.dout1 (dout_5_21),
	.dout1_valid (dout_valid_5_21)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_11 (
	.clk (clk),
	.addr0 (addr_5_22),
	.addr0_valid (addr_valid_5_22),
	.addr1 (addr_5_23),
	.addr1_valid (addr_valid_5_23),
	.dout0 (dout_5_22),
	.dout0_valid (dout_valid_5_22),
	.dout1 (dout_5_23),
	.dout1_valid (dout_valid_5_23)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_12 (
	.clk (clk),
	.addr0 (addr_5_24),
	.addr0_valid (addr_valid_5_24),
	.addr1 (addr_5_25),
	.addr1_valid (addr_valid_5_25),
	.dout0 (dout_5_24),
	.dout0_valid (dout_valid_5_24),
	.dout1 (dout_5_25),
	.dout1_valid (dout_valid_5_25)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_13 (
	.clk (clk),
	.addr0 (addr_5_26),
	.addr0_valid (addr_valid_5_26),
	.addr1 (addr_5_27),
	.addr1_valid (addr_valid_5_27),
	.dout0 (dout_5_26),
	.dout0_valid (dout_valid_5_26),
	.dout1 (dout_5_27),
	.dout1_valid (dout_valid_5_27)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_14 (
	.clk (clk),
	.addr0 (addr_5_28),
	.addr0_valid (addr_valid_5_28),
	.addr1 (addr_5_29),
	.addr1_valid (addr_valid_5_29),
	.dout0 (dout_5_28),
	.dout0_valid (dout_valid_5_28),
	.dout1 (dout_5_29),
	.dout1_valid (dout_valid_5_29)
);

hashtable #(
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./memory_init/bitmap5.mif")
)
hashtable_5_15 (
	.clk (clk),
	.addr0 (addr_5_30),
	.addr0_valid (addr_valid_5_30),
	.addr1 (addr_5_31),
	.addr1_valid (addr_valid_5_31),
	.dout0 (dout_5_30),
	.dout0_valid (dout_valid_5_30),
	.dout1 (dout_5_31),
	.dout1_valid (dout_valid_5_31)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_0 (
	.clk (clk),
	.addr0 (addr_6_0),
	.addr0_valid (addr_valid_6_0),
	.addr1 (addr_6_1),
	.addr1_valid (addr_valid_6_1),
	.dout0 (dout_6_0),
	.dout0_valid (dout_valid_6_0),
	.dout1 (dout_6_1),
	.dout1_valid (dout_valid_6_1)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_1 (
	.clk (clk),
	.addr0 (addr_6_2),
	.addr0_valid (addr_valid_6_2),
	.addr1 (addr_6_3),
	.addr1_valid (addr_valid_6_3),
	.dout0 (dout_6_2),
	.dout0_valid (dout_valid_6_2),
	.dout1 (dout_6_3),
	.dout1_valid (dout_valid_6_3)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_2 (
	.clk (clk),
	.addr0 (addr_6_4),
	.addr0_valid (addr_valid_6_4),
	.addr1 (addr_6_5),
	.addr1_valid (addr_valid_6_5),
	.dout0 (dout_6_4),
	.dout0_valid (dout_valid_6_4),
	.dout1 (dout_6_5),
	.dout1_valid (dout_valid_6_5)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_3 (
	.clk (clk),
	.addr0 (addr_6_6),
	.addr0_valid (addr_valid_6_6),
	.addr1 (addr_6_7),
	.addr1_valid (addr_valid_6_7),
	.dout0 (dout_6_6),
	.dout0_valid (dout_valid_6_6),
	.dout1 (dout_6_7),
	.dout1_valid (dout_valid_6_7)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_4 (
	.clk (clk),
	.addr0 (addr_6_8),
	.addr0_valid (addr_valid_6_8),
	.addr1 (addr_6_9),
	.addr1_valid (addr_valid_6_9),
	.dout0 (dout_6_8),
	.dout0_valid (dout_valid_6_8),
	.dout1 (dout_6_9),
	.dout1_valid (dout_valid_6_9)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_5 (
	.clk (clk),
	.addr0 (addr_6_10),
	.addr0_valid (addr_valid_6_10),
	.addr1 (addr_6_11),
	.addr1_valid (addr_valid_6_11),
	.dout0 (dout_6_10),
	.dout0_valid (dout_valid_6_10),
	.dout1 (dout_6_11),
	.dout1_valid (dout_valid_6_11)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_6 (
	.clk (clk),
	.addr0 (addr_6_12),
	.addr0_valid (addr_valid_6_12),
	.addr1 (addr_6_13),
	.addr1_valid (addr_valid_6_13),
	.dout0 (dout_6_12),
	.dout0_valid (dout_valid_6_12),
	.dout1 (dout_6_13),
	.dout1_valid (dout_valid_6_13)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_7 (
	.clk (clk),
	.addr0 (addr_6_14),
	.addr0_valid (addr_valid_6_14),
	.addr1 (addr_6_15),
	.addr1_valid (addr_valid_6_15),
	.dout0 (dout_6_14),
	.dout0_valid (dout_valid_6_14),
	.dout1 (dout_6_15),
	.dout1_valid (dout_valid_6_15)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_8 (
	.clk (clk),
	.addr0 (addr_6_16),
	.addr0_valid (addr_valid_6_16),
	.addr1 (addr_6_17),
	.addr1_valid (addr_valid_6_17),
	.dout0 (dout_6_16),
	.dout0_valid (dout_valid_6_16),
	.dout1 (dout_6_17),
	.dout1_valid (dout_valid_6_17)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_9 (
	.clk (clk),
	.addr0 (addr_6_18),
	.addr0_valid (addr_valid_6_18),
	.addr1 (addr_6_19),
	.addr1_valid (addr_valid_6_19),
	.dout0 (dout_6_18),
	.dout0_valid (dout_valid_6_18),
	.dout1 (dout_6_19),
	.dout1_valid (dout_valid_6_19)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_10 (
	.clk (clk),
	.addr0 (addr_6_20),
	.addr0_valid (addr_valid_6_20),
	.addr1 (addr_6_21),
	.addr1_valid (addr_valid_6_21),
	.dout0 (dout_6_20),
	.dout0_valid (dout_valid_6_20),
	.dout1 (dout_6_21),
	.dout1_valid (dout_valid_6_21)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_11 (
	.clk (clk),
	.addr0 (addr_6_22),
	.addr0_valid (addr_valid_6_22),
	.addr1 (addr_6_23),
	.addr1_valid (addr_valid_6_23),
	.dout0 (dout_6_22),
	.dout0_valid (dout_valid_6_22),
	.dout1 (dout_6_23),
	.dout1_valid (dout_valid_6_23)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_12 (
	.clk (clk),
	.addr0 (addr_6_24),
	.addr0_valid (addr_valid_6_24),
	.addr1 (addr_6_25),
	.addr1_valid (addr_valid_6_25),
	.dout0 (dout_6_24),
	.dout0_valid (dout_valid_6_24),
	.dout1 (dout_6_25),
	.dout1_valid (dout_valid_6_25)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_13 (
	.clk (clk),
	.addr0 (addr_6_26),
	.addr0_valid (addr_valid_6_26),
	.addr1 (addr_6_27),
	.addr1_valid (addr_valid_6_27),
	.dout0 (dout_6_26),
	.dout0_valid (dout_valid_6_26),
	.dout1 (dout_6_27),
	.dout1_valid (dout_valid_6_27)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_14 (
	.clk (clk),
	.addr0 (addr_6_28),
	.addr0_valid (addr_valid_6_28),
	.addr1 (addr_6_29),
	.addr1_valid (addr_valid_6_29),
	.dout0 (dout_6_28),
	.dout0_valid (dout_valid_6_28),
	.dout1 (dout_6_29),
	.dout1_valid (dout_valid_6_29)
);

hashtable #(
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./memory_init/bitmap6.mif")
)
hashtable_6_15 (
	.clk (clk),
	.addr0 (addr_6_30),
	.addr0_valid (addr_valid_6_30),
	.addr1 (addr_6_31),
	.addr1_valid (addr_valid_6_31),
	.dout0 (dout_6_30),
	.dout0_valid (dout_valid_6_30),
	.dout1 (dout_6_31),
	.dout1_valid (dout_valid_6_31)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_0 (
	.clk (clk),
	.addr0 (addr_7_0),
	.addr0_valid (addr_valid_7_0),
	.addr1 (addr_7_1),
	.addr1_valid (addr_valid_7_1),
	.dout0 (dout_7_0),
	.dout0_valid (dout_valid_7_0),
	.dout1 (dout_7_1),
	.dout1_valid (dout_valid_7_1)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_1 (
	.clk (clk),
	.addr0 (addr_7_2),
	.addr0_valid (addr_valid_7_2),
	.addr1 (addr_7_3),
	.addr1_valid (addr_valid_7_3),
	.dout0 (dout_7_2),
	.dout0_valid (dout_valid_7_2),
	.dout1 (dout_7_3),
	.dout1_valid (dout_valid_7_3)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_2 (
	.clk (clk),
	.addr0 (addr_7_4),
	.addr0_valid (addr_valid_7_4),
	.addr1 (addr_7_5),
	.addr1_valid (addr_valid_7_5),
	.dout0 (dout_7_4),
	.dout0_valid (dout_valid_7_4),
	.dout1 (dout_7_5),
	.dout1_valid (dout_valid_7_5)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_3 (
	.clk (clk),
	.addr0 (addr_7_6),
	.addr0_valid (addr_valid_7_6),
	.addr1 (addr_7_7),
	.addr1_valid (addr_valid_7_7),
	.dout0 (dout_7_6),
	.dout0_valid (dout_valid_7_6),
	.dout1 (dout_7_7),
	.dout1_valid (dout_valid_7_7)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_4 (
	.clk (clk),
	.addr0 (addr_7_8),
	.addr0_valid (addr_valid_7_8),
	.addr1 (addr_7_9),
	.addr1_valid (addr_valid_7_9),
	.dout0 (dout_7_8),
	.dout0_valid (dout_valid_7_8),
	.dout1 (dout_7_9),
	.dout1_valid (dout_valid_7_9)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_5 (
	.clk (clk),
	.addr0 (addr_7_10),
	.addr0_valid (addr_valid_7_10),
	.addr1 (addr_7_11),
	.addr1_valid (addr_valid_7_11),
	.dout0 (dout_7_10),
	.dout0_valid (dout_valid_7_10),
	.dout1 (dout_7_11),
	.dout1_valid (dout_valid_7_11)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_6 (
	.clk (clk),
	.addr0 (addr_7_12),
	.addr0_valid (addr_valid_7_12),
	.addr1 (addr_7_13),
	.addr1_valid (addr_valid_7_13),
	.dout0 (dout_7_12),
	.dout0_valid (dout_valid_7_12),
	.dout1 (dout_7_13),
	.dout1_valid (dout_valid_7_13)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_7 (
	.clk (clk),
	.addr0 (addr_7_14),
	.addr0_valid (addr_valid_7_14),
	.addr1 (addr_7_15),
	.addr1_valid (addr_valid_7_15),
	.dout0 (dout_7_14),
	.dout0_valid (dout_valid_7_14),
	.dout1 (dout_7_15),
	.dout1_valid (dout_valid_7_15)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_8 (
	.clk (clk),
	.addr0 (addr_7_16),
	.addr0_valid (addr_valid_7_16),
	.addr1 (addr_7_17),
	.addr1_valid (addr_valid_7_17),
	.dout0 (dout_7_16),
	.dout0_valid (dout_valid_7_16),
	.dout1 (dout_7_17),
	.dout1_valid (dout_valid_7_17)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_9 (
	.clk (clk),
	.addr0 (addr_7_18),
	.addr0_valid (addr_valid_7_18),
	.addr1 (addr_7_19),
	.addr1_valid (addr_valid_7_19),
	.dout0 (dout_7_18),
	.dout0_valid (dout_valid_7_18),
	.dout1 (dout_7_19),
	.dout1_valid (dout_valid_7_19)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_10 (
	.clk (clk),
	.addr0 (addr_7_20),
	.addr0_valid (addr_valid_7_20),
	.addr1 (addr_7_21),
	.addr1_valid (addr_valid_7_21),
	.dout0 (dout_7_20),
	.dout0_valid (dout_valid_7_20),
	.dout1 (dout_7_21),
	.dout1_valid (dout_valid_7_21)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_11 (
	.clk (clk),
	.addr0 (addr_7_22),
	.addr0_valid (addr_valid_7_22),
	.addr1 (addr_7_23),
	.addr1_valid (addr_valid_7_23),
	.dout0 (dout_7_22),
	.dout0_valid (dout_valid_7_22),
	.dout1 (dout_7_23),
	.dout1_valid (dout_valid_7_23)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_12 (
	.clk (clk),
	.addr0 (addr_7_24),
	.addr0_valid (addr_valid_7_24),
	.addr1 (addr_7_25),
	.addr1_valid (addr_valid_7_25),
	.dout0 (dout_7_24),
	.dout0_valid (dout_valid_7_24),
	.dout1 (dout_7_25),
	.dout1_valid (dout_valid_7_25)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_13 (
	.clk (clk),
	.addr0 (addr_7_26),
	.addr0_valid (addr_valid_7_26),
	.addr1 (addr_7_27),
	.addr1_valid (addr_valid_7_27),
	.dout0 (dout_7_26),
	.dout0_valid (dout_valid_7_26),
	.dout1 (dout_7_27),
	.dout1_valid (dout_valid_7_27)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_14 (
	.clk (clk),
	.addr0 (addr_7_28),
	.addr0_valid (addr_valid_7_28),
	.addr1 (addr_7_29),
	.addr1_valid (addr_valid_7_29),
	.dout0 (dout_7_28),
	.dout0_valid (dout_valid_7_28),
	.dout1 (dout_7_29),
	.dout1_valid (dout_valid_7_29)
);

hashtable #(
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./memory_init/bitmap7.mif")
)
hashtable_7_15 (
	.clk (clk),
	.addr0 (addr_7_30),
	.addr0_valid (addr_valid_7_30),
	.addr1 (addr_7_31),
	.addr1_valid (addr_valid_7_31),
	.dout0 (dout_7_30),
	.dout0_valid (dout_valid_7_30),
	.dout1 (dout_7_31),
	.dout1_valid (dout_valid_7_31)
);

endmodule
../../accel/pigasus_sme/rtl/struct_s.sv
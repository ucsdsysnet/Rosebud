`include "struct_s.sv"
module string_matcher (
    clk,
    rst,
    in_data,
    in_valid,
    in_sop,
    in_eop,
    in_empty,
    in_ready,
    in_meta_data,
    in_meta_valid,
    in_meta_ready,
    out_data,
    out_valid,
    out_almost_full,
    out_last,
    out_meta_data,
    out_meta_valid,
    out_meta_ready,
        // status register bus
    clk_status,
    status_addr,
    status_read,
    status_write,
    status_writedata,
    status_readdata,
    status_readdata_valid
);

input clk;
input rst;
input [255:0] in_data;
input in_valid;
input in_sop;
input in_eop;
input [4:0] in_empty;
output logic in_ready;
input metadata_t in_meta_data;
input in_meta_valid;
output logic in_meta_ready;
output metadata_t out_meta_data;
output logic out_meta_valid;
input logic out_meta_ready;
output logic [127:0] out_data;
output logic out_valid;
output logic out_last;
input out_almost_full;
// status register bus
input   logic          clk_status;
input   logic   [29:0] status_addr;
input   logic          status_read;
input   logic          status_write;
input   logic   [31:0] status_writedata;
output  logic   [31:0] status_readdata;
output  logic          status_readdata_valid;


logic [255:0] in_data_r1;
logic [255:0] in_data_r2;
logic         in_valid_r1;
logic         in_valid_r2;
logic         in_sop_r1;
logic         in_sop_r2;
logic         in_eop_r1;
logic         in_eop_r2;
logic [4:0]   in_empty_r1;
logic [4:0]   in_empty_r2;

metadata_t  internal_meta_data;
logic       internal_meta_valid;
logic       internal_meta_ready;

logic [RID_WIDTH-1:0] hash_out_0_0;
logic hash_out_valid_filter_0_0;
rule_s_t din_0_0;
rule_s_t din_0_0_r1;
rule_s_t din_0_0_r2;
logic din_valid_0_0;
logic din_valid_0_0_r1;
logic din_valid_0_0_r2;
logic [2:0] din_valid_0_0_r;
logic din_ready_0_0;
logic din_almost_full_0_0;
logic [RID_WIDTH-1:0] hash_out_0_1;
logic hash_out_valid_filter_0_1;
rule_s_t din_0_1;
rule_s_t din_0_1_r1;
rule_s_t din_0_1_r2;
logic din_valid_0_1;
logic din_valid_0_1_r1;
logic din_valid_0_1_r2;
logic [2:0] din_valid_0_1_r;
logic din_ready_0_1;
logic din_almost_full_0_1;
logic [RID_WIDTH-1:0] hash_out_0_2;
logic hash_out_valid_filter_0_2;
rule_s_t din_0_2;
rule_s_t din_0_2_r1;
rule_s_t din_0_2_r2;
logic din_valid_0_2;
logic din_valid_0_2_r1;
logic din_valid_0_2_r2;
logic [2:0] din_valid_0_2_r;
logic din_ready_0_2;
logic din_almost_full_0_2;
logic [RID_WIDTH-1:0] hash_out_0_3;
logic hash_out_valid_filter_0_3;
rule_s_t din_0_3;
rule_s_t din_0_3_r1;
rule_s_t din_0_3_r2;
logic din_valid_0_3;
logic din_valid_0_3_r1;
logic din_valid_0_3_r2;
logic [2:0] din_valid_0_3_r;
logic din_ready_0_3;
logic din_almost_full_0_3;
logic [RID_WIDTH-1:0] hash_out_0_4;
logic hash_out_valid_filter_0_4;
rule_s_t din_0_4;
rule_s_t din_0_4_r1;
rule_s_t din_0_4_r2;
logic din_valid_0_4;
logic din_valid_0_4_r1;
logic din_valid_0_4_r2;
logic [2:0] din_valid_0_4_r;
logic din_ready_0_4;
logic din_almost_full_0_4;
logic [RID_WIDTH-1:0] hash_out_0_5;
logic hash_out_valid_filter_0_5;
rule_s_t din_0_5;
rule_s_t din_0_5_r1;
rule_s_t din_0_5_r2;
logic din_valid_0_5;
logic din_valid_0_5_r1;
logic din_valid_0_5_r2;
logic [2:0] din_valid_0_5_r;
logic din_ready_0_5;
logic din_almost_full_0_5;
logic [RID_WIDTH-1:0] hash_out_0_6;
logic hash_out_valid_filter_0_6;
rule_s_t din_0_6;
rule_s_t din_0_6_r1;
rule_s_t din_0_6_r2;
logic din_valid_0_6;
logic din_valid_0_6_r1;
logic din_valid_0_6_r2;
logic [2:0] din_valid_0_6_r;
logic din_ready_0_6;
logic din_almost_full_0_6;
logic [RID_WIDTH-1:0] hash_out_0_7;
logic hash_out_valid_filter_0_7;
rule_s_t din_0_7;
rule_s_t din_0_7_r1;
rule_s_t din_0_7_r2;
logic din_valid_0_7;
logic din_valid_0_7_r1;
logic din_valid_0_7_r2;
logic [2:0] din_valid_0_7_r;
logic din_ready_0_7;
logic din_almost_full_0_7;
logic [RID_WIDTH-1:0] hash_out_0_8;
logic hash_out_valid_filter_0_8;
rule_s_t din_0_8;
rule_s_t din_0_8_r1;
rule_s_t din_0_8_r2;
logic din_valid_0_8;
logic din_valid_0_8_r1;
logic din_valid_0_8_r2;
logic [2:0] din_valid_0_8_r;
logic din_ready_0_8;
logic din_almost_full_0_8;
logic [RID_WIDTH-1:0] hash_out_0_9;
logic hash_out_valid_filter_0_9;
rule_s_t din_0_9;
rule_s_t din_0_9_r1;
rule_s_t din_0_9_r2;
logic din_valid_0_9;
logic din_valid_0_9_r1;
logic din_valid_0_9_r2;
logic [2:0] din_valid_0_9_r;
logic din_ready_0_9;
logic din_almost_full_0_9;
logic [RID_WIDTH-1:0] hash_out_0_10;
logic hash_out_valid_filter_0_10;
rule_s_t din_0_10;
rule_s_t din_0_10_r1;
rule_s_t din_0_10_r2;
logic din_valid_0_10;
logic din_valid_0_10_r1;
logic din_valid_0_10_r2;
logic [2:0] din_valid_0_10_r;
logic din_ready_0_10;
logic din_almost_full_0_10;
logic [RID_WIDTH-1:0] hash_out_0_11;
logic hash_out_valid_filter_0_11;
rule_s_t din_0_11;
rule_s_t din_0_11_r1;
rule_s_t din_0_11_r2;
logic din_valid_0_11;
logic din_valid_0_11_r1;
logic din_valid_0_11_r2;
logic [2:0] din_valid_0_11_r;
logic din_ready_0_11;
logic din_almost_full_0_11;
logic [RID_WIDTH-1:0] hash_out_0_12;
logic hash_out_valid_filter_0_12;
rule_s_t din_0_12;
rule_s_t din_0_12_r1;
rule_s_t din_0_12_r2;
logic din_valid_0_12;
logic din_valid_0_12_r1;
logic din_valid_0_12_r2;
logic [2:0] din_valid_0_12_r;
logic din_ready_0_12;
logic din_almost_full_0_12;
logic [RID_WIDTH-1:0] hash_out_0_13;
logic hash_out_valid_filter_0_13;
rule_s_t din_0_13;
rule_s_t din_0_13_r1;
rule_s_t din_0_13_r2;
logic din_valid_0_13;
logic din_valid_0_13_r1;
logic din_valid_0_13_r2;
logic [2:0] din_valid_0_13_r;
logic din_ready_0_13;
logic din_almost_full_0_13;
logic [RID_WIDTH-1:0] hash_out_0_14;
logic hash_out_valid_filter_0_14;
rule_s_t din_0_14;
rule_s_t din_0_14_r1;
rule_s_t din_0_14_r2;
logic din_valid_0_14;
logic din_valid_0_14_r1;
logic din_valid_0_14_r2;
logic [2:0] din_valid_0_14_r;
logic din_ready_0_14;
logic din_almost_full_0_14;
logic [RID_WIDTH-1:0] hash_out_0_15;
logic hash_out_valid_filter_0_15;
rule_s_t din_0_15;
rule_s_t din_0_15_r1;
rule_s_t din_0_15_r2;
logic din_valid_0_15;
logic din_valid_0_15_r1;
logic din_valid_0_15_r2;
logic [2:0] din_valid_0_15_r;
logic din_ready_0_15;
logic din_almost_full_0_15;
logic [RID_WIDTH-1:0] hash_out_0_16;
logic hash_out_valid_filter_0_16;
rule_s_t din_0_16;
rule_s_t din_0_16_r1;
rule_s_t din_0_16_r2;
logic din_valid_0_16;
logic din_valid_0_16_r1;
logic din_valid_0_16_r2;
logic [2:0] din_valid_0_16_r;
logic din_ready_0_16;
logic din_almost_full_0_16;
logic [RID_WIDTH-1:0] hash_out_0_17;
logic hash_out_valid_filter_0_17;
rule_s_t din_0_17;
rule_s_t din_0_17_r1;
rule_s_t din_0_17_r2;
logic din_valid_0_17;
logic din_valid_0_17_r1;
logic din_valid_0_17_r2;
logic [2:0] din_valid_0_17_r;
logic din_ready_0_17;
logic din_almost_full_0_17;
logic [RID_WIDTH-1:0] hash_out_0_18;
logic hash_out_valid_filter_0_18;
rule_s_t din_0_18;
rule_s_t din_0_18_r1;
rule_s_t din_0_18_r2;
logic din_valid_0_18;
logic din_valid_0_18_r1;
logic din_valid_0_18_r2;
logic [2:0] din_valid_0_18_r;
logic din_ready_0_18;
logic din_almost_full_0_18;
logic [RID_WIDTH-1:0] hash_out_0_19;
logic hash_out_valid_filter_0_19;
rule_s_t din_0_19;
rule_s_t din_0_19_r1;
rule_s_t din_0_19_r2;
logic din_valid_0_19;
logic din_valid_0_19_r1;
logic din_valid_0_19_r2;
logic [2:0] din_valid_0_19_r;
logic din_ready_0_19;
logic din_almost_full_0_19;
logic [RID_WIDTH-1:0] hash_out_0_20;
logic hash_out_valid_filter_0_20;
rule_s_t din_0_20;
rule_s_t din_0_20_r1;
rule_s_t din_0_20_r2;
logic din_valid_0_20;
logic din_valid_0_20_r1;
logic din_valid_0_20_r2;
logic [2:0] din_valid_0_20_r;
logic din_ready_0_20;
logic din_almost_full_0_20;
logic [RID_WIDTH-1:0] hash_out_0_21;
logic hash_out_valid_filter_0_21;
rule_s_t din_0_21;
rule_s_t din_0_21_r1;
rule_s_t din_0_21_r2;
logic din_valid_0_21;
logic din_valid_0_21_r1;
logic din_valid_0_21_r2;
logic [2:0] din_valid_0_21_r;
logic din_ready_0_21;
logic din_almost_full_0_21;
logic [RID_WIDTH-1:0] hash_out_0_22;
logic hash_out_valid_filter_0_22;
rule_s_t din_0_22;
rule_s_t din_0_22_r1;
rule_s_t din_0_22_r2;
logic din_valid_0_22;
logic din_valid_0_22_r1;
logic din_valid_0_22_r2;
logic [2:0] din_valid_0_22_r;
logic din_ready_0_22;
logic din_almost_full_0_22;
logic [RID_WIDTH-1:0] hash_out_0_23;
logic hash_out_valid_filter_0_23;
rule_s_t din_0_23;
rule_s_t din_0_23_r1;
rule_s_t din_0_23_r2;
logic din_valid_0_23;
logic din_valid_0_23_r1;
logic din_valid_0_23_r2;
logic [2:0] din_valid_0_23_r;
logic din_ready_0_23;
logic din_almost_full_0_23;
logic [RID_WIDTH-1:0] hash_out_0_24;
logic hash_out_valid_filter_0_24;
rule_s_t din_0_24;
rule_s_t din_0_24_r1;
rule_s_t din_0_24_r2;
logic din_valid_0_24;
logic din_valid_0_24_r1;
logic din_valid_0_24_r2;
logic [2:0] din_valid_0_24_r;
logic din_ready_0_24;
logic din_almost_full_0_24;
logic [RID_WIDTH-1:0] hash_out_0_25;
logic hash_out_valid_filter_0_25;
rule_s_t din_0_25;
rule_s_t din_0_25_r1;
rule_s_t din_0_25_r2;
logic din_valid_0_25;
logic din_valid_0_25_r1;
logic din_valid_0_25_r2;
logic [2:0] din_valid_0_25_r;
logic din_ready_0_25;
logic din_almost_full_0_25;
logic [RID_WIDTH-1:0] hash_out_0_26;
logic hash_out_valid_filter_0_26;
rule_s_t din_0_26;
rule_s_t din_0_26_r1;
rule_s_t din_0_26_r2;
logic din_valid_0_26;
logic din_valid_0_26_r1;
logic din_valid_0_26_r2;
logic [2:0] din_valid_0_26_r;
logic din_ready_0_26;
logic din_almost_full_0_26;
logic [RID_WIDTH-1:0] hash_out_0_27;
logic hash_out_valid_filter_0_27;
rule_s_t din_0_27;
rule_s_t din_0_27_r1;
rule_s_t din_0_27_r2;
logic din_valid_0_27;
logic din_valid_0_27_r1;
logic din_valid_0_27_r2;
logic [2:0] din_valid_0_27_r;
logic din_ready_0_27;
logic din_almost_full_0_27;
logic [RID_WIDTH-1:0] hash_out_0_28;
logic hash_out_valid_filter_0_28;
rule_s_t din_0_28;
rule_s_t din_0_28_r1;
rule_s_t din_0_28_r2;
logic din_valid_0_28;
logic din_valid_0_28_r1;
logic din_valid_0_28_r2;
logic [2:0] din_valid_0_28_r;
logic din_ready_0_28;
logic din_almost_full_0_28;
logic [RID_WIDTH-1:0] hash_out_0_29;
logic hash_out_valid_filter_0_29;
rule_s_t din_0_29;
rule_s_t din_0_29_r1;
rule_s_t din_0_29_r2;
logic din_valid_0_29;
logic din_valid_0_29_r1;
logic din_valid_0_29_r2;
logic [2:0] din_valid_0_29_r;
logic din_ready_0_29;
logic din_almost_full_0_29;
logic [RID_WIDTH-1:0] hash_out_0_30;
logic hash_out_valid_filter_0_30;
rule_s_t din_0_30;
rule_s_t din_0_30_r1;
rule_s_t din_0_30_r2;
logic din_valid_0_30;
logic din_valid_0_30_r1;
logic din_valid_0_30_r2;
logic [2:0] din_valid_0_30_r;
logic din_ready_0_30;
logic din_almost_full_0_30;
logic [RID_WIDTH-1:0] hash_out_0_31;
logic hash_out_valid_filter_0_31;
rule_s_t din_0_31;
rule_s_t din_0_31_r1;
rule_s_t din_0_31_r2;
logic din_valid_0_31;
logic din_valid_0_31_r1;
logic din_valid_0_31_r2;
logic [2:0] din_valid_0_31_r;
logic din_ready_0_31;
logic din_almost_full_0_31;
logic [RID_WIDTH-1:0] hash_out_1_0;
logic hash_out_valid_filter_1_0;
rule_s_t din_1_0;
rule_s_t din_1_0_r1;
rule_s_t din_1_0_r2;
logic din_valid_1_0;
logic din_valid_1_0_r1;
logic din_valid_1_0_r2;
logic [2:0] din_valid_1_0_r;
logic din_ready_1_0;
logic din_almost_full_1_0;
logic [RID_WIDTH-1:0] hash_out_1_1;
logic hash_out_valid_filter_1_1;
rule_s_t din_1_1;
rule_s_t din_1_1_r1;
rule_s_t din_1_1_r2;
logic din_valid_1_1;
logic din_valid_1_1_r1;
logic din_valid_1_1_r2;
logic [2:0] din_valid_1_1_r;
logic din_ready_1_1;
logic din_almost_full_1_1;
logic [RID_WIDTH-1:0] hash_out_1_2;
logic hash_out_valid_filter_1_2;
rule_s_t din_1_2;
rule_s_t din_1_2_r1;
rule_s_t din_1_2_r2;
logic din_valid_1_2;
logic din_valid_1_2_r1;
logic din_valid_1_2_r2;
logic [2:0] din_valid_1_2_r;
logic din_ready_1_2;
logic din_almost_full_1_2;
logic [RID_WIDTH-1:0] hash_out_1_3;
logic hash_out_valid_filter_1_3;
rule_s_t din_1_3;
rule_s_t din_1_3_r1;
rule_s_t din_1_3_r2;
logic din_valid_1_3;
logic din_valid_1_3_r1;
logic din_valid_1_3_r2;
logic [2:0] din_valid_1_3_r;
logic din_ready_1_3;
logic din_almost_full_1_3;
logic [RID_WIDTH-1:0] hash_out_1_4;
logic hash_out_valid_filter_1_4;
rule_s_t din_1_4;
rule_s_t din_1_4_r1;
rule_s_t din_1_4_r2;
logic din_valid_1_4;
logic din_valid_1_4_r1;
logic din_valid_1_4_r2;
logic [2:0] din_valid_1_4_r;
logic din_ready_1_4;
logic din_almost_full_1_4;
logic [RID_WIDTH-1:0] hash_out_1_5;
logic hash_out_valid_filter_1_5;
rule_s_t din_1_5;
rule_s_t din_1_5_r1;
rule_s_t din_1_5_r2;
logic din_valid_1_5;
logic din_valid_1_5_r1;
logic din_valid_1_5_r2;
logic [2:0] din_valid_1_5_r;
logic din_ready_1_5;
logic din_almost_full_1_5;
logic [RID_WIDTH-1:0] hash_out_1_6;
logic hash_out_valid_filter_1_6;
rule_s_t din_1_6;
rule_s_t din_1_6_r1;
rule_s_t din_1_6_r2;
logic din_valid_1_6;
logic din_valid_1_6_r1;
logic din_valid_1_6_r2;
logic [2:0] din_valid_1_6_r;
logic din_ready_1_6;
logic din_almost_full_1_6;
logic [RID_WIDTH-1:0] hash_out_1_7;
logic hash_out_valid_filter_1_7;
rule_s_t din_1_7;
rule_s_t din_1_7_r1;
rule_s_t din_1_7_r2;
logic din_valid_1_7;
logic din_valid_1_7_r1;
logic din_valid_1_7_r2;
logic [2:0] din_valid_1_7_r;
logic din_ready_1_7;
logic din_almost_full_1_7;
logic [RID_WIDTH-1:0] hash_out_1_8;
logic hash_out_valid_filter_1_8;
rule_s_t din_1_8;
rule_s_t din_1_8_r1;
rule_s_t din_1_8_r2;
logic din_valid_1_8;
logic din_valid_1_8_r1;
logic din_valid_1_8_r2;
logic [2:0] din_valid_1_8_r;
logic din_ready_1_8;
logic din_almost_full_1_8;
logic [RID_WIDTH-1:0] hash_out_1_9;
logic hash_out_valid_filter_1_9;
rule_s_t din_1_9;
rule_s_t din_1_9_r1;
rule_s_t din_1_9_r2;
logic din_valid_1_9;
logic din_valid_1_9_r1;
logic din_valid_1_9_r2;
logic [2:0] din_valid_1_9_r;
logic din_ready_1_9;
logic din_almost_full_1_9;
logic [RID_WIDTH-1:0] hash_out_1_10;
logic hash_out_valid_filter_1_10;
rule_s_t din_1_10;
rule_s_t din_1_10_r1;
rule_s_t din_1_10_r2;
logic din_valid_1_10;
logic din_valid_1_10_r1;
logic din_valid_1_10_r2;
logic [2:0] din_valid_1_10_r;
logic din_ready_1_10;
logic din_almost_full_1_10;
logic [RID_WIDTH-1:0] hash_out_1_11;
logic hash_out_valid_filter_1_11;
rule_s_t din_1_11;
rule_s_t din_1_11_r1;
rule_s_t din_1_11_r2;
logic din_valid_1_11;
logic din_valid_1_11_r1;
logic din_valid_1_11_r2;
logic [2:0] din_valid_1_11_r;
logic din_ready_1_11;
logic din_almost_full_1_11;
logic [RID_WIDTH-1:0] hash_out_1_12;
logic hash_out_valid_filter_1_12;
rule_s_t din_1_12;
rule_s_t din_1_12_r1;
rule_s_t din_1_12_r2;
logic din_valid_1_12;
logic din_valid_1_12_r1;
logic din_valid_1_12_r2;
logic [2:0] din_valid_1_12_r;
logic din_ready_1_12;
logic din_almost_full_1_12;
logic [RID_WIDTH-1:0] hash_out_1_13;
logic hash_out_valid_filter_1_13;
rule_s_t din_1_13;
rule_s_t din_1_13_r1;
rule_s_t din_1_13_r2;
logic din_valid_1_13;
logic din_valid_1_13_r1;
logic din_valid_1_13_r2;
logic [2:0] din_valid_1_13_r;
logic din_ready_1_13;
logic din_almost_full_1_13;
logic [RID_WIDTH-1:0] hash_out_1_14;
logic hash_out_valid_filter_1_14;
rule_s_t din_1_14;
rule_s_t din_1_14_r1;
rule_s_t din_1_14_r2;
logic din_valid_1_14;
logic din_valid_1_14_r1;
logic din_valid_1_14_r2;
logic [2:0] din_valid_1_14_r;
logic din_ready_1_14;
logic din_almost_full_1_14;
logic [RID_WIDTH-1:0] hash_out_1_15;
logic hash_out_valid_filter_1_15;
rule_s_t din_1_15;
rule_s_t din_1_15_r1;
rule_s_t din_1_15_r2;
logic din_valid_1_15;
logic din_valid_1_15_r1;
logic din_valid_1_15_r2;
logic [2:0] din_valid_1_15_r;
logic din_ready_1_15;
logic din_almost_full_1_15;
logic [RID_WIDTH-1:0] hash_out_1_16;
logic hash_out_valid_filter_1_16;
rule_s_t din_1_16;
rule_s_t din_1_16_r1;
rule_s_t din_1_16_r2;
logic din_valid_1_16;
logic din_valid_1_16_r1;
logic din_valid_1_16_r2;
logic [2:0] din_valid_1_16_r;
logic din_ready_1_16;
logic din_almost_full_1_16;
logic [RID_WIDTH-1:0] hash_out_1_17;
logic hash_out_valid_filter_1_17;
rule_s_t din_1_17;
rule_s_t din_1_17_r1;
rule_s_t din_1_17_r2;
logic din_valid_1_17;
logic din_valid_1_17_r1;
logic din_valid_1_17_r2;
logic [2:0] din_valid_1_17_r;
logic din_ready_1_17;
logic din_almost_full_1_17;
logic [RID_WIDTH-1:0] hash_out_1_18;
logic hash_out_valid_filter_1_18;
rule_s_t din_1_18;
rule_s_t din_1_18_r1;
rule_s_t din_1_18_r2;
logic din_valid_1_18;
logic din_valid_1_18_r1;
logic din_valid_1_18_r2;
logic [2:0] din_valid_1_18_r;
logic din_ready_1_18;
logic din_almost_full_1_18;
logic [RID_WIDTH-1:0] hash_out_1_19;
logic hash_out_valid_filter_1_19;
rule_s_t din_1_19;
rule_s_t din_1_19_r1;
rule_s_t din_1_19_r2;
logic din_valid_1_19;
logic din_valid_1_19_r1;
logic din_valid_1_19_r2;
logic [2:0] din_valid_1_19_r;
logic din_ready_1_19;
logic din_almost_full_1_19;
logic [RID_WIDTH-1:0] hash_out_1_20;
logic hash_out_valid_filter_1_20;
rule_s_t din_1_20;
rule_s_t din_1_20_r1;
rule_s_t din_1_20_r2;
logic din_valid_1_20;
logic din_valid_1_20_r1;
logic din_valid_1_20_r2;
logic [2:0] din_valid_1_20_r;
logic din_ready_1_20;
logic din_almost_full_1_20;
logic [RID_WIDTH-1:0] hash_out_1_21;
logic hash_out_valid_filter_1_21;
rule_s_t din_1_21;
rule_s_t din_1_21_r1;
rule_s_t din_1_21_r2;
logic din_valid_1_21;
logic din_valid_1_21_r1;
logic din_valid_1_21_r2;
logic [2:0] din_valid_1_21_r;
logic din_ready_1_21;
logic din_almost_full_1_21;
logic [RID_WIDTH-1:0] hash_out_1_22;
logic hash_out_valid_filter_1_22;
rule_s_t din_1_22;
rule_s_t din_1_22_r1;
rule_s_t din_1_22_r2;
logic din_valid_1_22;
logic din_valid_1_22_r1;
logic din_valid_1_22_r2;
logic [2:0] din_valid_1_22_r;
logic din_ready_1_22;
logic din_almost_full_1_22;
logic [RID_WIDTH-1:0] hash_out_1_23;
logic hash_out_valid_filter_1_23;
rule_s_t din_1_23;
rule_s_t din_1_23_r1;
rule_s_t din_1_23_r2;
logic din_valid_1_23;
logic din_valid_1_23_r1;
logic din_valid_1_23_r2;
logic [2:0] din_valid_1_23_r;
logic din_ready_1_23;
logic din_almost_full_1_23;
logic [RID_WIDTH-1:0] hash_out_1_24;
logic hash_out_valid_filter_1_24;
rule_s_t din_1_24;
rule_s_t din_1_24_r1;
rule_s_t din_1_24_r2;
logic din_valid_1_24;
logic din_valid_1_24_r1;
logic din_valid_1_24_r2;
logic [2:0] din_valid_1_24_r;
logic din_ready_1_24;
logic din_almost_full_1_24;
logic [RID_WIDTH-1:0] hash_out_1_25;
logic hash_out_valid_filter_1_25;
rule_s_t din_1_25;
rule_s_t din_1_25_r1;
rule_s_t din_1_25_r2;
logic din_valid_1_25;
logic din_valid_1_25_r1;
logic din_valid_1_25_r2;
logic [2:0] din_valid_1_25_r;
logic din_ready_1_25;
logic din_almost_full_1_25;
logic [RID_WIDTH-1:0] hash_out_1_26;
logic hash_out_valid_filter_1_26;
rule_s_t din_1_26;
rule_s_t din_1_26_r1;
rule_s_t din_1_26_r2;
logic din_valid_1_26;
logic din_valid_1_26_r1;
logic din_valid_1_26_r2;
logic [2:0] din_valid_1_26_r;
logic din_ready_1_26;
logic din_almost_full_1_26;
logic [RID_WIDTH-1:0] hash_out_1_27;
logic hash_out_valid_filter_1_27;
rule_s_t din_1_27;
rule_s_t din_1_27_r1;
rule_s_t din_1_27_r2;
logic din_valid_1_27;
logic din_valid_1_27_r1;
logic din_valid_1_27_r2;
logic [2:0] din_valid_1_27_r;
logic din_ready_1_27;
logic din_almost_full_1_27;
logic [RID_WIDTH-1:0] hash_out_1_28;
logic hash_out_valid_filter_1_28;
rule_s_t din_1_28;
rule_s_t din_1_28_r1;
rule_s_t din_1_28_r2;
logic din_valid_1_28;
logic din_valid_1_28_r1;
logic din_valid_1_28_r2;
logic [2:0] din_valid_1_28_r;
logic din_ready_1_28;
logic din_almost_full_1_28;
logic [RID_WIDTH-1:0] hash_out_1_29;
logic hash_out_valid_filter_1_29;
rule_s_t din_1_29;
rule_s_t din_1_29_r1;
rule_s_t din_1_29_r2;
logic din_valid_1_29;
logic din_valid_1_29_r1;
logic din_valid_1_29_r2;
logic [2:0] din_valid_1_29_r;
logic din_ready_1_29;
logic din_almost_full_1_29;
logic [RID_WIDTH-1:0] hash_out_1_30;
logic hash_out_valid_filter_1_30;
rule_s_t din_1_30;
rule_s_t din_1_30_r1;
rule_s_t din_1_30_r2;
logic din_valid_1_30;
logic din_valid_1_30_r1;
logic din_valid_1_30_r2;
logic [2:0] din_valid_1_30_r;
logic din_ready_1_30;
logic din_almost_full_1_30;
logic [RID_WIDTH-1:0] hash_out_1_31;
logic hash_out_valid_filter_1_31;
rule_s_t din_1_31;
rule_s_t din_1_31_r1;
rule_s_t din_1_31_r2;
logic din_valid_1_31;
logic din_valid_1_31_r1;
logic din_valid_1_31_r2;
logic [2:0] din_valid_1_31_r;
logic din_ready_1_31;
logic din_almost_full_1_31;
logic [RID_WIDTH-1:0] hash_out_2_0;
logic hash_out_valid_filter_2_0;
rule_s_t din_2_0;
rule_s_t din_2_0_r1;
rule_s_t din_2_0_r2;
logic din_valid_2_0;
logic din_valid_2_0_r1;
logic din_valid_2_0_r2;
logic [2:0] din_valid_2_0_r;
logic din_ready_2_0;
logic din_almost_full_2_0;
logic [RID_WIDTH-1:0] hash_out_2_1;
logic hash_out_valid_filter_2_1;
rule_s_t din_2_1;
rule_s_t din_2_1_r1;
rule_s_t din_2_1_r2;
logic din_valid_2_1;
logic din_valid_2_1_r1;
logic din_valid_2_1_r2;
logic [2:0] din_valid_2_1_r;
logic din_ready_2_1;
logic din_almost_full_2_1;
logic [RID_WIDTH-1:0] hash_out_2_2;
logic hash_out_valid_filter_2_2;
rule_s_t din_2_2;
rule_s_t din_2_2_r1;
rule_s_t din_2_2_r2;
logic din_valid_2_2;
logic din_valid_2_2_r1;
logic din_valid_2_2_r2;
logic [2:0] din_valid_2_2_r;
logic din_ready_2_2;
logic din_almost_full_2_2;
logic [RID_WIDTH-1:0] hash_out_2_3;
logic hash_out_valid_filter_2_3;
rule_s_t din_2_3;
rule_s_t din_2_3_r1;
rule_s_t din_2_3_r2;
logic din_valid_2_3;
logic din_valid_2_3_r1;
logic din_valid_2_3_r2;
logic [2:0] din_valid_2_3_r;
logic din_ready_2_3;
logic din_almost_full_2_3;
logic [RID_WIDTH-1:0] hash_out_2_4;
logic hash_out_valid_filter_2_4;
rule_s_t din_2_4;
rule_s_t din_2_4_r1;
rule_s_t din_2_4_r2;
logic din_valid_2_4;
logic din_valid_2_4_r1;
logic din_valid_2_4_r2;
logic [2:0] din_valid_2_4_r;
logic din_ready_2_4;
logic din_almost_full_2_4;
logic [RID_WIDTH-1:0] hash_out_2_5;
logic hash_out_valid_filter_2_5;
rule_s_t din_2_5;
rule_s_t din_2_5_r1;
rule_s_t din_2_5_r2;
logic din_valid_2_5;
logic din_valid_2_5_r1;
logic din_valid_2_5_r2;
logic [2:0] din_valid_2_5_r;
logic din_ready_2_5;
logic din_almost_full_2_5;
logic [RID_WIDTH-1:0] hash_out_2_6;
logic hash_out_valid_filter_2_6;
rule_s_t din_2_6;
rule_s_t din_2_6_r1;
rule_s_t din_2_6_r2;
logic din_valid_2_6;
logic din_valid_2_6_r1;
logic din_valid_2_6_r2;
logic [2:0] din_valid_2_6_r;
logic din_ready_2_6;
logic din_almost_full_2_6;
logic [RID_WIDTH-1:0] hash_out_2_7;
logic hash_out_valid_filter_2_7;
rule_s_t din_2_7;
rule_s_t din_2_7_r1;
rule_s_t din_2_7_r2;
logic din_valid_2_7;
logic din_valid_2_7_r1;
logic din_valid_2_7_r2;
logic [2:0] din_valid_2_7_r;
logic din_ready_2_7;
logic din_almost_full_2_7;
logic [RID_WIDTH-1:0] hash_out_2_8;
logic hash_out_valid_filter_2_8;
rule_s_t din_2_8;
rule_s_t din_2_8_r1;
rule_s_t din_2_8_r2;
logic din_valid_2_8;
logic din_valid_2_8_r1;
logic din_valid_2_8_r2;
logic [2:0] din_valid_2_8_r;
logic din_ready_2_8;
logic din_almost_full_2_8;
logic [RID_WIDTH-1:0] hash_out_2_9;
logic hash_out_valid_filter_2_9;
rule_s_t din_2_9;
rule_s_t din_2_9_r1;
rule_s_t din_2_9_r2;
logic din_valid_2_9;
logic din_valid_2_9_r1;
logic din_valid_2_9_r2;
logic [2:0] din_valid_2_9_r;
logic din_ready_2_9;
logic din_almost_full_2_9;
logic [RID_WIDTH-1:0] hash_out_2_10;
logic hash_out_valid_filter_2_10;
rule_s_t din_2_10;
rule_s_t din_2_10_r1;
rule_s_t din_2_10_r2;
logic din_valid_2_10;
logic din_valid_2_10_r1;
logic din_valid_2_10_r2;
logic [2:0] din_valid_2_10_r;
logic din_ready_2_10;
logic din_almost_full_2_10;
logic [RID_WIDTH-1:0] hash_out_2_11;
logic hash_out_valid_filter_2_11;
rule_s_t din_2_11;
rule_s_t din_2_11_r1;
rule_s_t din_2_11_r2;
logic din_valid_2_11;
logic din_valid_2_11_r1;
logic din_valid_2_11_r2;
logic [2:0] din_valid_2_11_r;
logic din_ready_2_11;
logic din_almost_full_2_11;
logic [RID_WIDTH-1:0] hash_out_2_12;
logic hash_out_valid_filter_2_12;
rule_s_t din_2_12;
rule_s_t din_2_12_r1;
rule_s_t din_2_12_r2;
logic din_valid_2_12;
logic din_valid_2_12_r1;
logic din_valid_2_12_r2;
logic [2:0] din_valid_2_12_r;
logic din_ready_2_12;
logic din_almost_full_2_12;
logic [RID_WIDTH-1:0] hash_out_2_13;
logic hash_out_valid_filter_2_13;
rule_s_t din_2_13;
rule_s_t din_2_13_r1;
rule_s_t din_2_13_r2;
logic din_valid_2_13;
logic din_valid_2_13_r1;
logic din_valid_2_13_r2;
logic [2:0] din_valid_2_13_r;
logic din_ready_2_13;
logic din_almost_full_2_13;
logic [RID_WIDTH-1:0] hash_out_2_14;
logic hash_out_valid_filter_2_14;
rule_s_t din_2_14;
rule_s_t din_2_14_r1;
rule_s_t din_2_14_r2;
logic din_valid_2_14;
logic din_valid_2_14_r1;
logic din_valid_2_14_r2;
logic [2:0] din_valid_2_14_r;
logic din_ready_2_14;
logic din_almost_full_2_14;
logic [RID_WIDTH-1:0] hash_out_2_15;
logic hash_out_valid_filter_2_15;
rule_s_t din_2_15;
rule_s_t din_2_15_r1;
rule_s_t din_2_15_r2;
logic din_valid_2_15;
logic din_valid_2_15_r1;
logic din_valid_2_15_r2;
logic [2:0] din_valid_2_15_r;
logic din_ready_2_15;
logic din_almost_full_2_15;
logic [RID_WIDTH-1:0] hash_out_2_16;
logic hash_out_valid_filter_2_16;
rule_s_t din_2_16;
rule_s_t din_2_16_r1;
rule_s_t din_2_16_r2;
logic din_valid_2_16;
logic din_valid_2_16_r1;
logic din_valid_2_16_r2;
logic [2:0] din_valid_2_16_r;
logic din_ready_2_16;
logic din_almost_full_2_16;
logic [RID_WIDTH-1:0] hash_out_2_17;
logic hash_out_valid_filter_2_17;
rule_s_t din_2_17;
rule_s_t din_2_17_r1;
rule_s_t din_2_17_r2;
logic din_valid_2_17;
logic din_valid_2_17_r1;
logic din_valid_2_17_r2;
logic [2:0] din_valid_2_17_r;
logic din_ready_2_17;
logic din_almost_full_2_17;
logic [RID_WIDTH-1:0] hash_out_2_18;
logic hash_out_valid_filter_2_18;
rule_s_t din_2_18;
rule_s_t din_2_18_r1;
rule_s_t din_2_18_r2;
logic din_valid_2_18;
logic din_valid_2_18_r1;
logic din_valid_2_18_r2;
logic [2:0] din_valid_2_18_r;
logic din_ready_2_18;
logic din_almost_full_2_18;
logic [RID_WIDTH-1:0] hash_out_2_19;
logic hash_out_valid_filter_2_19;
rule_s_t din_2_19;
rule_s_t din_2_19_r1;
rule_s_t din_2_19_r2;
logic din_valid_2_19;
logic din_valid_2_19_r1;
logic din_valid_2_19_r2;
logic [2:0] din_valid_2_19_r;
logic din_ready_2_19;
logic din_almost_full_2_19;
logic [RID_WIDTH-1:0] hash_out_2_20;
logic hash_out_valid_filter_2_20;
rule_s_t din_2_20;
rule_s_t din_2_20_r1;
rule_s_t din_2_20_r2;
logic din_valid_2_20;
logic din_valid_2_20_r1;
logic din_valid_2_20_r2;
logic [2:0] din_valid_2_20_r;
logic din_ready_2_20;
logic din_almost_full_2_20;
logic [RID_WIDTH-1:0] hash_out_2_21;
logic hash_out_valid_filter_2_21;
rule_s_t din_2_21;
rule_s_t din_2_21_r1;
rule_s_t din_2_21_r2;
logic din_valid_2_21;
logic din_valid_2_21_r1;
logic din_valid_2_21_r2;
logic [2:0] din_valid_2_21_r;
logic din_ready_2_21;
logic din_almost_full_2_21;
logic [RID_WIDTH-1:0] hash_out_2_22;
logic hash_out_valid_filter_2_22;
rule_s_t din_2_22;
rule_s_t din_2_22_r1;
rule_s_t din_2_22_r2;
logic din_valid_2_22;
logic din_valid_2_22_r1;
logic din_valid_2_22_r2;
logic [2:0] din_valid_2_22_r;
logic din_ready_2_22;
logic din_almost_full_2_22;
logic [RID_WIDTH-1:0] hash_out_2_23;
logic hash_out_valid_filter_2_23;
rule_s_t din_2_23;
rule_s_t din_2_23_r1;
rule_s_t din_2_23_r2;
logic din_valid_2_23;
logic din_valid_2_23_r1;
logic din_valid_2_23_r2;
logic [2:0] din_valid_2_23_r;
logic din_ready_2_23;
logic din_almost_full_2_23;
logic [RID_WIDTH-1:0] hash_out_2_24;
logic hash_out_valid_filter_2_24;
rule_s_t din_2_24;
rule_s_t din_2_24_r1;
rule_s_t din_2_24_r2;
logic din_valid_2_24;
logic din_valid_2_24_r1;
logic din_valid_2_24_r2;
logic [2:0] din_valid_2_24_r;
logic din_ready_2_24;
logic din_almost_full_2_24;
logic [RID_WIDTH-1:0] hash_out_2_25;
logic hash_out_valid_filter_2_25;
rule_s_t din_2_25;
rule_s_t din_2_25_r1;
rule_s_t din_2_25_r2;
logic din_valid_2_25;
logic din_valid_2_25_r1;
logic din_valid_2_25_r2;
logic [2:0] din_valid_2_25_r;
logic din_ready_2_25;
logic din_almost_full_2_25;
logic [RID_WIDTH-1:0] hash_out_2_26;
logic hash_out_valid_filter_2_26;
rule_s_t din_2_26;
rule_s_t din_2_26_r1;
rule_s_t din_2_26_r2;
logic din_valid_2_26;
logic din_valid_2_26_r1;
logic din_valid_2_26_r2;
logic [2:0] din_valid_2_26_r;
logic din_ready_2_26;
logic din_almost_full_2_26;
logic [RID_WIDTH-1:0] hash_out_2_27;
logic hash_out_valid_filter_2_27;
rule_s_t din_2_27;
rule_s_t din_2_27_r1;
rule_s_t din_2_27_r2;
logic din_valid_2_27;
logic din_valid_2_27_r1;
logic din_valid_2_27_r2;
logic [2:0] din_valid_2_27_r;
logic din_ready_2_27;
logic din_almost_full_2_27;
logic [RID_WIDTH-1:0] hash_out_2_28;
logic hash_out_valid_filter_2_28;
rule_s_t din_2_28;
rule_s_t din_2_28_r1;
rule_s_t din_2_28_r2;
logic din_valid_2_28;
logic din_valid_2_28_r1;
logic din_valid_2_28_r2;
logic [2:0] din_valid_2_28_r;
logic din_ready_2_28;
logic din_almost_full_2_28;
logic [RID_WIDTH-1:0] hash_out_2_29;
logic hash_out_valid_filter_2_29;
rule_s_t din_2_29;
rule_s_t din_2_29_r1;
rule_s_t din_2_29_r2;
logic din_valid_2_29;
logic din_valid_2_29_r1;
logic din_valid_2_29_r2;
logic [2:0] din_valid_2_29_r;
logic din_ready_2_29;
logic din_almost_full_2_29;
logic [RID_WIDTH-1:0] hash_out_2_30;
logic hash_out_valid_filter_2_30;
rule_s_t din_2_30;
rule_s_t din_2_30_r1;
rule_s_t din_2_30_r2;
logic din_valid_2_30;
logic din_valid_2_30_r1;
logic din_valid_2_30_r2;
logic [2:0] din_valid_2_30_r;
logic din_ready_2_30;
logic din_almost_full_2_30;
logic [RID_WIDTH-1:0] hash_out_2_31;
logic hash_out_valid_filter_2_31;
rule_s_t din_2_31;
rule_s_t din_2_31_r1;
rule_s_t din_2_31_r2;
logic din_valid_2_31;
logic din_valid_2_31_r1;
logic din_valid_2_31_r2;
logic [2:0] din_valid_2_31_r;
logic din_ready_2_31;
logic din_almost_full_2_31;
logic [RID_WIDTH-1:0] hash_out_3_0;
logic hash_out_valid_filter_3_0;
rule_s_t din_3_0;
rule_s_t din_3_0_r1;
rule_s_t din_3_0_r2;
logic din_valid_3_0;
logic din_valid_3_0_r1;
logic din_valid_3_0_r2;
logic [2:0] din_valid_3_0_r;
logic din_ready_3_0;
logic din_almost_full_3_0;
logic [RID_WIDTH-1:0] hash_out_3_1;
logic hash_out_valid_filter_3_1;
rule_s_t din_3_1;
rule_s_t din_3_1_r1;
rule_s_t din_3_1_r2;
logic din_valid_3_1;
logic din_valid_3_1_r1;
logic din_valid_3_1_r2;
logic [2:0] din_valid_3_1_r;
logic din_ready_3_1;
logic din_almost_full_3_1;
logic [RID_WIDTH-1:0] hash_out_3_2;
logic hash_out_valid_filter_3_2;
rule_s_t din_3_2;
rule_s_t din_3_2_r1;
rule_s_t din_3_2_r2;
logic din_valid_3_2;
logic din_valid_3_2_r1;
logic din_valid_3_2_r2;
logic [2:0] din_valid_3_2_r;
logic din_ready_3_2;
logic din_almost_full_3_2;
logic [RID_WIDTH-1:0] hash_out_3_3;
logic hash_out_valid_filter_3_3;
rule_s_t din_3_3;
rule_s_t din_3_3_r1;
rule_s_t din_3_3_r2;
logic din_valid_3_3;
logic din_valid_3_3_r1;
logic din_valid_3_3_r2;
logic [2:0] din_valid_3_3_r;
logic din_ready_3_3;
logic din_almost_full_3_3;
logic [RID_WIDTH-1:0] hash_out_3_4;
logic hash_out_valid_filter_3_4;
rule_s_t din_3_4;
rule_s_t din_3_4_r1;
rule_s_t din_3_4_r2;
logic din_valid_3_4;
logic din_valid_3_4_r1;
logic din_valid_3_4_r2;
logic [2:0] din_valid_3_4_r;
logic din_ready_3_4;
logic din_almost_full_3_4;
logic [RID_WIDTH-1:0] hash_out_3_5;
logic hash_out_valid_filter_3_5;
rule_s_t din_3_5;
rule_s_t din_3_5_r1;
rule_s_t din_3_5_r2;
logic din_valid_3_5;
logic din_valid_3_5_r1;
logic din_valid_3_5_r2;
logic [2:0] din_valid_3_5_r;
logic din_ready_3_5;
logic din_almost_full_3_5;
logic [RID_WIDTH-1:0] hash_out_3_6;
logic hash_out_valid_filter_3_6;
rule_s_t din_3_6;
rule_s_t din_3_6_r1;
rule_s_t din_3_6_r2;
logic din_valid_3_6;
logic din_valid_3_6_r1;
logic din_valid_3_6_r2;
logic [2:0] din_valid_3_6_r;
logic din_ready_3_6;
logic din_almost_full_3_6;
logic [RID_WIDTH-1:0] hash_out_3_7;
logic hash_out_valid_filter_3_7;
rule_s_t din_3_7;
rule_s_t din_3_7_r1;
rule_s_t din_3_7_r2;
logic din_valid_3_7;
logic din_valid_3_7_r1;
logic din_valid_3_7_r2;
logic [2:0] din_valid_3_7_r;
logic din_ready_3_7;
logic din_almost_full_3_7;
logic [RID_WIDTH-1:0] hash_out_3_8;
logic hash_out_valid_filter_3_8;
rule_s_t din_3_8;
rule_s_t din_3_8_r1;
rule_s_t din_3_8_r2;
logic din_valid_3_8;
logic din_valid_3_8_r1;
logic din_valid_3_8_r2;
logic [2:0] din_valid_3_8_r;
logic din_ready_3_8;
logic din_almost_full_3_8;
logic [RID_WIDTH-1:0] hash_out_3_9;
logic hash_out_valid_filter_3_9;
rule_s_t din_3_9;
rule_s_t din_3_9_r1;
rule_s_t din_3_9_r2;
logic din_valid_3_9;
logic din_valid_3_9_r1;
logic din_valid_3_9_r2;
logic [2:0] din_valid_3_9_r;
logic din_ready_3_9;
logic din_almost_full_3_9;
logic [RID_WIDTH-1:0] hash_out_3_10;
logic hash_out_valid_filter_3_10;
rule_s_t din_3_10;
rule_s_t din_3_10_r1;
rule_s_t din_3_10_r2;
logic din_valid_3_10;
logic din_valid_3_10_r1;
logic din_valid_3_10_r2;
logic [2:0] din_valid_3_10_r;
logic din_ready_3_10;
logic din_almost_full_3_10;
logic [RID_WIDTH-1:0] hash_out_3_11;
logic hash_out_valid_filter_3_11;
rule_s_t din_3_11;
rule_s_t din_3_11_r1;
rule_s_t din_3_11_r2;
logic din_valid_3_11;
logic din_valid_3_11_r1;
logic din_valid_3_11_r2;
logic [2:0] din_valid_3_11_r;
logic din_ready_3_11;
logic din_almost_full_3_11;
logic [RID_WIDTH-1:0] hash_out_3_12;
logic hash_out_valid_filter_3_12;
rule_s_t din_3_12;
rule_s_t din_3_12_r1;
rule_s_t din_3_12_r2;
logic din_valid_3_12;
logic din_valid_3_12_r1;
logic din_valid_3_12_r2;
logic [2:0] din_valid_3_12_r;
logic din_ready_3_12;
logic din_almost_full_3_12;
logic [RID_WIDTH-1:0] hash_out_3_13;
logic hash_out_valid_filter_3_13;
rule_s_t din_3_13;
rule_s_t din_3_13_r1;
rule_s_t din_3_13_r2;
logic din_valid_3_13;
logic din_valid_3_13_r1;
logic din_valid_3_13_r2;
logic [2:0] din_valid_3_13_r;
logic din_ready_3_13;
logic din_almost_full_3_13;
logic [RID_WIDTH-1:0] hash_out_3_14;
logic hash_out_valid_filter_3_14;
rule_s_t din_3_14;
rule_s_t din_3_14_r1;
rule_s_t din_3_14_r2;
logic din_valid_3_14;
logic din_valid_3_14_r1;
logic din_valid_3_14_r2;
logic [2:0] din_valid_3_14_r;
logic din_ready_3_14;
logic din_almost_full_3_14;
logic [RID_WIDTH-1:0] hash_out_3_15;
logic hash_out_valid_filter_3_15;
rule_s_t din_3_15;
rule_s_t din_3_15_r1;
rule_s_t din_3_15_r2;
logic din_valid_3_15;
logic din_valid_3_15_r1;
logic din_valid_3_15_r2;
logic [2:0] din_valid_3_15_r;
logic din_ready_3_15;
logic din_almost_full_3_15;
logic [RID_WIDTH-1:0] hash_out_3_16;
logic hash_out_valid_filter_3_16;
rule_s_t din_3_16;
rule_s_t din_3_16_r1;
rule_s_t din_3_16_r2;
logic din_valid_3_16;
logic din_valid_3_16_r1;
logic din_valid_3_16_r2;
logic [2:0] din_valid_3_16_r;
logic din_ready_3_16;
logic din_almost_full_3_16;
logic [RID_WIDTH-1:0] hash_out_3_17;
logic hash_out_valid_filter_3_17;
rule_s_t din_3_17;
rule_s_t din_3_17_r1;
rule_s_t din_3_17_r2;
logic din_valid_3_17;
logic din_valid_3_17_r1;
logic din_valid_3_17_r2;
logic [2:0] din_valid_3_17_r;
logic din_ready_3_17;
logic din_almost_full_3_17;
logic [RID_WIDTH-1:0] hash_out_3_18;
logic hash_out_valid_filter_3_18;
rule_s_t din_3_18;
rule_s_t din_3_18_r1;
rule_s_t din_3_18_r2;
logic din_valid_3_18;
logic din_valid_3_18_r1;
logic din_valid_3_18_r2;
logic [2:0] din_valid_3_18_r;
logic din_ready_3_18;
logic din_almost_full_3_18;
logic [RID_WIDTH-1:0] hash_out_3_19;
logic hash_out_valid_filter_3_19;
rule_s_t din_3_19;
rule_s_t din_3_19_r1;
rule_s_t din_3_19_r2;
logic din_valid_3_19;
logic din_valid_3_19_r1;
logic din_valid_3_19_r2;
logic [2:0] din_valid_3_19_r;
logic din_ready_3_19;
logic din_almost_full_3_19;
logic [RID_WIDTH-1:0] hash_out_3_20;
logic hash_out_valid_filter_3_20;
rule_s_t din_3_20;
rule_s_t din_3_20_r1;
rule_s_t din_3_20_r2;
logic din_valid_3_20;
logic din_valid_3_20_r1;
logic din_valid_3_20_r2;
logic [2:0] din_valid_3_20_r;
logic din_ready_3_20;
logic din_almost_full_3_20;
logic [RID_WIDTH-1:0] hash_out_3_21;
logic hash_out_valid_filter_3_21;
rule_s_t din_3_21;
rule_s_t din_3_21_r1;
rule_s_t din_3_21_r2;
logic din_valid_3_21;
logic din_valid_3_21_r1;
logic din_valid_3_21_r2;
logic [2:0] din_valid_3_21_r;
logic din_ready_3_21;
logic din_almost_full_3_21;
logic [RID_WIDTH-1:0] hash_out_3_22;
logic hash_out_valid_filter_3_22;
rule_s_t din_3_22;
rule_s_t din_3_22_r1;
rule_s_t din_3_22_r2;
logic din_valid_3_22;
logic din_valid_3_22_r1;
logic din_valid_3_22_r2;
logic [2:0] din_valid_3_22_r;
logic din_ready_3_22;
logic din_almost_full_3_22;
logic [RID_WIDTH-1:0] hash_out_3_23;
logic hash_out_valid_filter_3_23;
rule_s_t din_3_23;
rule_s_t din_3_23_r1;
rule_s_t din_3_23_r2;
logic din_valid_3_23;
logic din_valid_3_23_r1;
logic din_valid_3_23_r2;
logic [2:0] din_valid_3_23_r;
logic din_ready_3_23;
logic din_almost_full_3_23;
logic [RID_WIDTH-1:0] hash_out_3_24;
logic hash_out_valid_filter_3_24;
rule_s_t din_3_24;
rule_s_t din_3_24_r1;
rule_s_t din_3_24_r2;
logic din_valid_3_24;
logic din_valid_3_24_r1;
logic din_valid_3_24_r2;
logic [2:0] din_valid_3_24_r;
logic din_ready_3_24;
logic din_almost_full_3_24;
logic [RID_WIDTH-1:0] hash_out_3_25;
logic hash_out_valid_filter_3_25;
rule_s_t din_3_25;
rule_s_t din_3_25_r1;
rule_s_t din_3_25_r2;
logic din_valid_3_25;
logic din_valid_3_25_r1;
logic din_valid_3_25_r2;
logic [2:0] din_valid_3_25_r;
logic din_ready_3_25;
logic din_almost_full_3_25;
logic [RID_WIDTH-1:0] hash_out_3_26;
logic hash_out_valid_filter_3_26;
rule_s_t din_3_26;
rule_s_t din_3_26_r1;
rule_s_t din_3_26_r2;
logic din_valid_3_26;
logic din_valid_3_26_r1;
logic din_valid_3_26_r2;
logic [2:0] din_valid_3_26_r;
logic din_ready_3_26;
logic din_almost_full_3_26;
logic [RID_WIDTH-1:0] hash_out_3_27;
logic hash_out_valid_filter_3_27;
rule_s_t din_3_27;
rule_s_t din_3_27_r1;
rule_s_t din_3_27_r2;
logic din_valid_3_27;
logic din_valid_3_27_r1;
logic din_valid_3_27_r2;
logic [2:0] din_valid_3_27_r;
logic din_ready_3_27;
logic din_almost_full_3_27;
logic [RID_WIDTH-1:0] hash_out_3_28;
logic hash_out_valid_filter_3_28;
rule_s_t din_3_28;
rule_s_t din_3_28_r1;
rule_s_t din_3_28_r2;
logic din_valid_3_28;
logic din_valid_3_28_r1;
logic din_valid_3_28_r2;
logic [2:0] din_valid_3_28_r;
logic din_ready_3_28;
logic din_almost_full_3_28;
logic [RID_WIDTH-1:0] hash_out_3_29;
logic hash_out_valid_filter_3_29;
rule_s_t din_3_29;
rule_s_t din_3_29_r1;
rule_s_t din_3_29_r2;
logic din_valid_3_29;
logic din_valid_3_29_r1;
logic din_valid_3_29_r2;
logic [2:0] din_valid_3_29_r;
logic din_ready_3_29;
logic din_almost_full_3_29;
logic [RID_WIDTH-1:0] hash_out_3_30;
logic hash_out_valid_filter_3_30;
rule_s_t din_3_30;
rule_s_t din_3_30_r1;
rule_s_t din_3_30_r2;
logic din_valid_3_30;
logic din_valid_3_30_r1;
logic din_valid_3_30_r2;
logic [2:0] din_valid_3_30_r;
logic din_ready_3_30;
logic din_almost_full_3_30;
logic [RID_WIDTH-1:0] hash_out_3_31;
logic hash_out_valid_filter_3_31;
rule_s_t din_3_31;
rule_s_t din_3_31_r1;
rule_s_t din_3_31_r2;
logic din_valid_3_31;
logic din_valid_3_31_r1;
logic din_valid_3_31_r2;
logic [2:0] din_valid_3_31_r;
logic din_ready_3_31;
logic din_almost_full_3_31;
logic [RID_WIDTH-1:0] hash_out_4_0;
logic hash_out_valid_filter_4_0;
rule_s_t din_4_0;
rule_s_t din_4_0_r1;
rule_s_t din_4_0_r2;
logic din_valid_4_0;
logic din_valid_4_0_r1;
logic din_valid_4_0_r2;
logic [2:0] din_valid_4_0_r;
logic din_ready_4_0;
logic din_almost_full_4_0;
logic [RID_WIDTH-1:0] hash_out_4_1;
logic hash_out_valid_filter_4_1;
rule_s_t din_4_1;
rule_s_t din_4_1_r1;
rule_s_t din_4_1_r2;
logic din_valid_4_1;
logic din_valid_4_1_r1;
logic din_valid_4_1_r2;
logic [2:0] din_valid_4_1_r;
logic din_ready_4_1;
logic din_almost_full_4_1;
logic [RID_WIDTH-1:0] hash_out_4_2;
logic hash_out_valid_filter_4_2;
rule_s_t din_4_2;
rule_s_t din_4_2_r1;
rule_s_t din_4_2_r2;
logic din_valid_4_2;
logic din_valid_4_2_r1;
logic din_valid_4_2_r2;
logic [2:0] din_valid_4_2_r;
logic din_ready_4_2;
logic din_almost_full_4_2;
logic [RID_WIDTH-1:0] hash_out_4_3;
logic hash_out_valid_filter_4_3;
rule_s_t din_4_3;
rule_s_t din_4_3_r1;
rule_s_t din_4_3_r2;
logic din_valid_4_3;
logic din_valid_4_3_r1;
logic din_valid_4_3_r2;
logic [2:0] din_valid_4_3_r;
logic din_ready_4_3;
logic din_almost_full_4_3;
logic [RID_WIDTH-1:0] hash_out_4_4;
logic hash_out_valid_filter_4_4;
rule_s_t din_4_4;
rule_s_t din_4_4_r1;
rule_s_t din_4_4_r2;
logic din_valid_4_4;
logic din_valid_4_4_r1;
logic din_valid_4_4_r2;
logic [2:0] din_valid_4_4_r;
logic din_ready_4_4;
logic din_almost_full_4_4;
logic [RID_WIDTH-1:0] hash_out_4_5;
logic hash_out_valid_filter_4_5;
rule_s_t din_4_5;
rule_s_t din_4_5_r1;
rule_s_t din_4_5_r2;
logic din_valid_4_5;
logic din_valid_4_5_r1;
logic din_valid_4_5_r2;
logic [2:0] din_valid_4_5_r;
logic din_ready_4_5;
logic din_almost_full_4_5;
logic [RID_WIDTH-1:0] hash_out_4_6;
logic hash_out_valid_filter_4_6;
rule_s_t din_4_6;
rule_s_t din_4_6_r1;
rule_s_t din_4_6_r2;
logic din_valid_4_6;
logic din_valid_4_6_r1;
logic din_valid_4_6_r2;
logic [2:0] din_valid_4_6_r;
logic din_ready_4_6;
logic din_almost_full_4_6;
logic [RID_WIDTH-1:0] hash_out_4_7;
logic hash_out_valid_filter_4_7;
rule_s_t din_4_7;
rule_s_t din_4_7_r1;
rule_s_t din_4_7_r2;
logic din_valid_4_7;
logic din_valid_4_7_r1;
logic din_valid_4_7_r2;
logic [2:0] din_valid_4_7_r;
logic din_ready_4_7;
logic din_almost_full_4_7;
logic [RID_WIDTH-1:0] hash_out_4_8;
logic hash_out_valid_filter_4_8;
rule_s_t din_4_8;
rule_s_t din_4_8_r1;
rule_s_t din_4_8_r2;
logic din_valid_4_8;
logic din_valid_4_8_r1;
logic din_valid_4_8_r2;
logic [2:0] din_valid_4_8_r;
logic din_ready_4_8;
logic din_almost_full_4_8;
logic [RID_WIDTH-1:0] hash_out_4_9;
logic hash_out_valid_filter_4_9;
rule_s_t din_4_9;
rule_s_t din_4_9_r1;
rule_s_t din_4_9_r2;
logic din_valid_4_9;
logic din_valid_4_9_r1;
logic din_valid_4_9_r2;
logic [2:0] din_valid_4_9_r;
logic din_ready_4_9;
logic din_almost_full_4_9;
logic [RID_WIDTH-1:0] hash_out_4_10;
logic hash_out_valid_filter_4_10;
rule_s_t din_4_10;
rule_s_t din_4_10_r1;
rule_s_t din_4_10_r2;
logic din_valid_4_10;
logic din_valid_4_10_r1;
logic din_valid_4_10_r2;
logic [2:0] din_valid_4_10_r;
logic din_ready_4_10;
logic din_almost_full_4_10;
logic [RID_WIDTH-1:0] hash_out_4_11;
logic hash_out_valid_filter_4_11;
rule_s_t din_4_11;
rule_s_t din_4_11_r1;
rule_s_t din_4_11_r2;
logic din_valid_4_11;
logic din_valid_4_11_r1;
logic din_valid_4_11_r2;
logic [2:0] din_valid_4_11_r;
logic din_ready_4_11;
logic din_almost_full_4_11;
logic [RID_WIDTH-1:0] hash_out_4_12;
logic hash_out_valid_filter_4_12;
rule_s_t din_4_12;
rule_s_t din_4_12_r1;
rule_s_t din_4_12_r2;
logic din_valid_4_12;
logic din_valid_4_12_r1;
logic din_valid_4_12_r2;
logic [2:0] din_valid_4_12_r;
logic din_ready_4_12;
logic din_almost_full_4_12;
logic [RID_WIDTH-1:0] hash_out_4_13;
logic hash_out_valid_filter_4_13;
rule_s_t din_4_13;
rule_s_t din_4_13_r1;
rule_s_t din_4_13_r2;
logic din_valid_4_13;
logic din_valid_4_13_r1;
logic din_valid_4_13_r2;
logic [2:0] din_valid_4_13_r;
logic din_ready_4_13;
logic din_almost_full_4_13;
logic [RID_WIDTH-1:0] hash_out_4_14;
logic hash_out_valid_filter_4_14;
rule_s_t din_4_14;
rule_s_t din_4_14_r1;
rule_s_t din_4_14_r2;
logic din_valid_4_14;
logic din_valid_4_14_r1;
logic din_valid_4_14_r2;
logic [2:0] din_valid_4_14_r;
logic din_ready_4_14;
logic din_almost_full_4_14;
logic [RID_WIDTH-1:0] hash_out_4_15;
logic hash_out_valid_filter_4_15;
rule_s_t din_4_15;
rule_s_t din_4_15_r1;
rule_s_t din_4_15_r2;
logic din_valid_4_15;
logic din_valid_4_15_r1;
logic din_valid_4_15_r2;
logic [2:0] din_valid_4_15_r;
logic din_ready_4_15;
logic din_almost_full_4_15;
logic [RID_WIDTH-1:0] hash_out_4_16;
logic hash_out_valid_filter_4_16;
rule_s_t din_4_16;
rule_s_t din_4_16_r1;
rule_s_t din_4_16_r2;
logic din_valid_4_16;
logic din_valid_4_16_r1;
logic din_valid_4_16_r2;
logic [2:0] din_valid_4_16_r;
logic din_ready_4_16;
logic din_almost_full_4_16;
logic [RID_WIDTH-1:0] hash_out_4_17;
logic hash_out_valid_filter_4_17;
rule_s_t din_4_17;
rule_s_t din_4_17_r1;
rule_s_t din_4_17_r2;
logic din_valid_4_17;
logic din_valid_4_17_r1;
logic din_valid_4_17_r2;
logic [2:0] din_valid_4_17_r;
logic din_ready_4_17;
logic din_almost_full_4_17;
logic [RID_WIDTH-1:0] hash_out_4_18;
logic hash_out_valid_filter_4_18;
rule_s_t din_4_18;
rule_s_t din_4_18_r1;
rule_s_t din_4_18_r2;
logic din_valid_4_18;
logic din_valid_4_18_r1;
logic din_valid_4_18_r2;
logic [2:0] din_valid_4_18_r;
logic din_ready_4_18;
logic din_almost_full_4_18;
logic [RID_WIDTH-1:0] hash_out_4_19;
logic hash_out_valid_filter_4_19;
rule_s_t din_4_19;
rule_s_t din_4_19_r1;
rule_s_t din_4_19_r2;
logic din_valid_4_19;
logic din_valid_4_19_r1;
logic din_valid_4_19_r2;
logic [2:0] din_valid_4_19_r;
logic din_ready_4_19;
logic din_almost_full_4_19;
logic [RID_WIDTH-1:0] hash_out_4_20;
logic hash_out_valid_filter_4_20;
rule_s_t din_4_20;
rule_s_t din_4_20_r1;
rule_s_t din_4_20_r2;
logic din_valid_4_20;
logic din_valid_4_20_r1;
logic din_valid_4_20_r2;
logic [2:0] din_valid_4_20_r;
logic din_ready_4_20;
logic din_almost_full_4_20;
logic [RID_WIDTH-1:0] hash_out_4_21;
logic hash_out_valid_filter_4_21;
rule_s_t din_4_21;
rule_s_t din_4_21_r1;
rule_s_t din_4_21_r2;
logic din_valid_4_21;
logic din_valid_4_21_r1;
logic din_valid_4_21_r2;
logic [2:0] din_valid_4_21_r;
logic din_ready_4_21;
logic din_almost_full_4_21;
logic [RID_WIDTH-1:0] hash_out_4_22;
logic hash_out_valid_filter_4_22;
rule_s_t din_4_22;
rule_s_t din_4_22_r1;
rule_s_t din_4_22_r2;
logic din_valid_4_22;
logic din_valid_4_22_r1;
logic din_valid_4_22_r2;
logic [2:0] din_valid_4_22_r;
logic din_ready_4_22;
logic din_almost_full_4_22;
logic [RID_WIDTH-1:0] hash_out_4_23;
logic hash_out_valid_filter_4_23;
rule_s_t din_4_23;
rule_s_t din_4_23_r1;
rule_s_t din_4_23_r2;
logic din_valid_4_23;
logic din_valid_4_23_r1;
logic din_valid_4_23_r2;
logic [2:0] din_valid_4_23_r;
logic din_ready_4_23;
logic din_almost_full_4_23;
logic [RID_WIDTH-1:0] hash_out_4_24;
logic hash_out_valid_filter_4_24;
rule_s_t din_4_24;
rule_s_t din_4_24_r1;
rule_s_t din_4_24_r2;
logic din_valid_4_24;
logic din_valid_4_24_r1;
logic din_valid_4_24_r2;
logic [2:0] din_valid_4_24_r;
logic din_ready_4_24;
logic din_almost_full_4_24;
logic [RID_WIDTH-1:0] hash_out_4_25;
logic hash_out_valid_filter_4_25;
rule_s_t din_4_25;
rule_s_t din_4_25_r1;
rule_s_t din_4_25_r2;
logic din_valid_4_25;
logic din_valid_4_25_r1;
logic din_valid_4_25_r2;
logic [2:0] din_valid_4_25_r;
logic din_ready_4_25;
logic din_almost_full_4_25;
logic [RID_WIDTH-1:0] hash_out_4_26;
logic hash_out_valid_filter_4_26;
rule_s_t din_4_26;
rule_s_t din_4_26_r1;
rule_s_t din_4_26_r2;
logic din_valid_4_26;
logic din_valid_4_26_r1;
logic din_valid_4_26_r2;
logic [2:0] din_valid_4_26_r;
logic din_ready_4_26;
logic din_almost_full_4_26;
logic [RID_WIDTH-1:0] hash_out_4_27;
logic hash_out_valid_filter_4_27;
rule_s_t din_4_27;
rule_s_t din_4_27_r1;
rule_s_t din_4_27_r2;
logic din_valid_4_27;
logic din_valid_4_27_r1;
logic din_valid_4_27_r2;
logic [2:0] din_valid_4_27_r;
logic din_ready_4_27;
logic din_almost_full_4_27;
logic [RID_WIDTH-1:0] hash_out_4_28;
logic hash_out_valid_filter_4_28;
rule_s_t din_4_28;
rule_s_t din_4_28_r1;
rule_s_t din_4_28_r2;
logic din_valid_4_28;
logic din_valid_4_28_r1;
logic din_valid_4_28_r2;
logic [2:0] din_valid_4_28_r;
logic din_ready_4_28;
logic din_almost_full_4_28;
logic [RID_WIDTH-1:0] hash_out_4_29;
logic hash_out_valid_filter_4_29;
rule_s_t din_4_29;
rule_s_t din_4_29_r1;
rule_s_t din_4_29_r2;
logic din_valid_4_29;
logic din_valid_4_29_r1;
logic din_valid_4_29_r2;
logic [2:0] din_valid_4_29_r;
logic din_ready_4_29;
logic din_almost_full_4_29;
logic [RID_WIDTH-1:0] hash_out_4_30;
logic hash_out_valid_filter_4_30;
rule_s_t din_4_30;
rule_s_t din_4_30_r1;
rule_s_t din_4_30_r2;
logic din_valid_4_30;
logic din_valid_4_30_r1;
logic din_valid_4_30_r2;
logic [2:0] din_valid_4_30_r;
logic din_ready_4_30;
logic din_almost_full_4_30;
logic [RID_WIDTH-1:0] hash_out_4_31;
logic hash_out_valid_filter_4_31;
rule_s_t din_4_31;
rule_s_t din_4_31_r1;
rule_s_t din_4_31_r2;
logic din_valid_4_31;
logic din_valid_4_31_r1;
logic din_valid_4_31_r2;
logic [2:0] din_valid_4_31_r;
logic din_ready_4_31;
logic din_almost_full_4_31;
logic [RID_WIDTH-1:0] hash_out_5_0;
logic hash_out_valid_filter_5_0;
rule_s_t din_5_0;
rule_s_t din_5_0_r1;
rule_s_t din_5_0_r2;
logic din_valid_5_0;
logic din_valid_5_0_r1;
logic din_valid_5_0_r2;
logic [2:0] din_valid_5_0_r;
logic din_ready_5_0;
logic din_almost_full_5_0;
logic [RID_WIDTH-1:0] hash_out_5_1;
logic hash_out_valid_filter_5_1;
rule_s_t din_5_1;
rule_s_t din_5_1_r1;
rule_s_t din_5_1_r2;
logic din_valid_5_1;
logic din_valid_5_1_r1;
logic din_valid_5_1_r2;
logic [2:0] din_valid_5_1_r;
logic din_ready_5_1;
logic din_almost_full_5_1;
logic [RID_WIDTH-1:0] hash_out_5_2;
logic hash_out_valid_filter_5_2;
rule_s_t din_5_2;
rule_s_t din_5_2_r1;
rule_s_t din_5_2_r2;
logic din_valid_5_2;
logic din_valid_5_2_r1;
logic din_valid_5_2_r2;
logic [2:0] din_valid_5_2_r;
logic din_ready_5_2;
logic din_almost_full_5_2;
logic [RID_WIDTH-1:0] hash_out_5_3;
logic hash_out_valid_filter_5_3;
rule_s_t din_5_3;
rule_s_t din_5_3_r1;
rule_s_t din_5_3_r2;
logic din_valid_5_3;
logic din_valid_5_3_r1;
logic din_valid_5_3_r2;
logic [2:0] din_valid_5_3_r;
logic din_ready_5_3;
logic din_almost_full_5_3;
logic [RID_WIDTH-1:0] hash_out_5_4;
logic hash_out_valid_filter_5_4;
rule_s_t din_5_4;
rule_s_t din_5_4_r1;
rule_s_t din_5_4_r2;
logic din_valid_5_4;
logic din_valid_5_4_r1;
logic din_valid_5_4_r2;
logic [2:0] din_valid_5_4_r;
logic din_ready_5_4;
logic din_almost_full_5_4;
logic [RID_WIDTH-1:0] hash_out_5_5;
logic hash_out_valid_filter_5_5;
rule_s_t din_5_5;
rule_s_t din_5_5_r1;
rule_s_t din_5_5_r2;
logic din_valid_5_5;
logic din_valid_5_5_r1;
logic din_valid_5_5_r2;
logic [2:0] din_valid_5_5_r;
logic din_ready_5_5;
logic din_almost_full_5_5;
logic [RID_WIDTH-1:0] hash_out_5_6;
logic hash_out_valid_filter_5_6;
rule_s_t din_5_6;
rule_s_t din_5_6_r1;
rule_s_t din_5_6_r2;
logic din_valid_5_6;
logic din_valid_5_6_r1;
logic din_valid_5_6_r2;
logic [2:0] din_valid_5_6_r;
logic din_ready_5_6;
logic din_almost_full_5_6;
logic [RID_WIDTH-1:0] hash_out_5_7;
logic hash_out_valid_filter_5_7;
rule_s_t din_5_7;
rule_s_t din_5_7_r1;
rule_s_t din_5_7_r2;
logic din_valid_5_7;
logic din_valid_5_7_r1;
logic din_valid_5_7_r2;
logic [2:0] din_valid_5_7_r;
logic din_ready_5_7;
logic din_almost_full_5_7;
logic [RID_WIDTH-1:0] hash_out_5_8;
logic hash_out_valid_filter_5_8;
rule_s_t din_5_8;
rule_s_t din_5_8_r1;
rule_s_t din_5_8_r2;
logic din_valid_5_8;
logic din_valid_5_8_r1;
logic din_valid_5_8_r2;
logic [2:0] din_valid_5_8_r;
logic din_ready_5_8;
logic din_almost_full_5_8;
logic [RID_WIDTH-1:0] hash_out_5_9;
logic hash_out_valid_filter_5_9;
rule_s_t din_5_9;
rule_s_t din_5_9_r1;
rule_s_t din_5_9_r2;
logic din_valid_5_9;
logic din_valid_5_9_r1;
logic din_valid_5_9_r2;
logic [2:0] din_valid_5_9_r;
logic din_ready_5_9;
logic din_almost_full_5_9;
logic [RID_WIDTH-1:0] hash_out_5_10;
logic hash_out_valid_filter_5_10;
rule_s_t din_5_10;
rule_s_t din_5_10_r1;
rule_s_t din_5_10_r2;
logic din_valid_5_10;
logic din_valid_5_10_r1;
logic din_valid_5_10_r2;
logic [2:0] din_valid_5_10_r;
logic din_ready_5_10;
logic din_almost_full_5_10;
logic [RID_WIDTH-1:0] hash_out_5_11;
logic hash_out_valid_filter_5_11;
rule_s_t din_5_11;
rule_s_t din_5_11_r1;
rule_s_t din_5_11_r2;
logic din_valid_5_11;
logic din_valid_5_11_r1;
logic din_valid_5_11_r2;
logic [2:0] din_valid_5_11_r;
logic din_ready_5_11;
logic din_almost_full_5_11;
logic [RID_WIDTH-1:0] hash_out_5_12;
logic hash_out_valid_filter_5_12;
rule_s_t din_5_12;
rule_s_t din_5_12_r1;
rule_s_t din_5_12_r2;
logic din_valid_5_12;
logic din_valid_5_12_r1;
logic din_valid_5_12_r2;
logic [2:0] din_valid_5_12_r;
logic din_ready_5_12;
logic din_almost_full_5_12;
logic [RID_WIDTH-1:0] hash_out_5_13;
logic hash_out_valid_filter_5_13;
rule_s_t din_5_13;
rule_s_t din_5_13_r1;
rule_s_t din_5_13_r2;
logic din_valid_5_13;
logic din_valid_5_13_r1;
logic din_valid_5_13_r2;
logic [2:0] din_valid_5_13_r;
logic din_ready_5_13;
logic din_almost_full_5_13;
logic [RID_WIDTH-1:0] hash_out_5_14;
logic hash_out_valid_filter_5_14;
rule_s_t din_5_14;
rule_s_t din_5_14_r1;
rule_s_t din_5_14_r2;
logic din_valid_5_14;
logic din_valid_5_14_r1;
logic din_valid_5_14_r2;
logic [2:0] din_valid_5_14_r;
logic din_ready_5_14;
logic din_almost_full_5_14;
logic [RID_WIDTH-1:0] hash_out_5_15;
logic hash_out_valid_filter_5_15;
rule_s_t din_5_15;
rule_s_t din_5_15_r1;
rule_s_t din_5_15_r2;
logic din_valid_5_15;
logic din_valid_5_15_r1;
logic din_valid_5_15_r2;
logic [2:0] din_valid_5_15_r;
logic din_ready_5_15;
logic din_almost_full_5_15;
logic [RID_WIDTH-1:0] hash_out_5_16;
logic hash_out_valid_filter_5_16;
rule_s_t din_5_16;
rule_s_t din_5_16_r1;
rule_s_t din_5_16_r2;
logic din_valid_5_16;
logic din_valid_5_16_r1;
logic din_valid_5_16_r2;
logic [2:0] din_valid_5_16_r;
logic din_ready_5_16;
logic din_almost_full_5_16;
logic [RID_WIDTH-1:0] hash_out_5_17;
logic hash_out_valid_filter_5_17;
rule_s_t din_5_17;
rule_s_t din_5_17_r1;
rule_s_t din_5_17_r2;
logic din_valid_5_17;
logic din_valid_5_17_r1;
logic din_valid_5_17_r2;
logic [2:0] din_valid_5_17_r;
logic din_ready_5_17;
logic din_almost_full_5_17;
logic [RID_WIDTH-1:0] hash_out_5_18;
logic hash_out_valid_filter_5_18;
rule_s_t din_5_18;
rule_s_t din_5_18_r1;
rule_s_t din_5_18_r2;
logic din_valid_5_18;
logic din_valid_5_18_r1;
logic din_valid_5_18_r2;
logic [2:0] din_valid_5_18_r;
logic din_ready_5_18;
logic din_almost_full_5_18;
logic [RID_WIDTH-1:0] hash_out_5_19;
logic hash_out_valid_filter_5_19;
rule_s_t din_5_19;
rule_s_t din_5_19_r1;
rule_s_t din_5_19_r2;
logic din_valid_5_19;
logic din_valid_5_19_r1;
logic din_valid_5_19_r2;
logic [2:0] din_valid_5_19_r;
logic din_ready_5_19;
logic din_almost_full_5_19;
logic [RID_WIDTH-1:0] hash_out_5_20;
logic hash_out_valid_filter_5_20;
rule_s_t din_5_20;
rule_s_t din_5_20_r1;
rule_s_t din_5_20_r2;
logic din_valid_5_20;
logic din_valid_5_20_r1;
logic din_valid_5_20_r2;
logic [2:0] din_valid_5_20_r;
logic din_ready_5_20;
logic din_almost_full_5_20;
logic [RID_WIDTH-1:0] hash_out_5_21;
logic hash_out_valid_filter_5_21;
rule_s_t din_5_21;
rule_s_t din_5_21_r1;
rule_s_t din_5_21_r2;
logic din_valid_5_21;
logic din_valid_5_21_r1;
logic din_valid_5_21_r2;
logic [2:0] din_valid_5_21_r;
logic din_ready_5_21;
logic din_almost_full_5_21;
logic [RID_WIDTH-1:0] hash_out_5_22;
logic hash_out_valid_filter_5_22;
rule_s_t din_5_22;
rule_s_t din_5_22_r1;
rule_s_t din_5_22_r2;
logic din_valid_5_22;
logic din_valid_5_22_r1;
logic din_valid_5_22_r2;
logic [2:0] din_valid_5_22_r;
logic din_ready_5_22;
logic din_almost_full_5_22;
logic [RID_WIDTH-1:0] hash_out_5_23;
logic hash_out_valid_filter_5_23;
rule_s_t din_5_23;
rule_s_t din_5_23_r1;
rule_s_t din_5_23_r2;
logic din_valid_5_23;
logic din_valid_5_23_r1;
logic din_valid_5_23_r2;
logic [2:0] din_valid_5_23_r;
logic din_ready_5_23;
logic din_almost_full_5_23;
logic [RID_WIDTH-1:0] hash_out_5_24;
logic hash_out_valid_filter_5_24;
rule_s_t din_5_24;
rule_s_t din_5_24_r1;
rule_s_t din_5_24_r2;
logic din_valid_5_24;
logic din_valid_5_24_r1;
logic din_valid_5_24_r2;
logic [2:0] din_valid_5_24_r;
logic din_ready_5_24;
logic din_almost_full_5_24;
logic [RID_WIDTH-1:0] hash_out_5_25;
logic hash_out_valid_filter_5_25;
rule_s_t din_5_25;
rule_s_t din_5_25_r1;
rule_s_t din_5_25_r2;
logic din_valid_5_25;
logic din_valid_5_25_r1;
logic din_valid_5_25_r2;
logic [2:0] din_valid_5_25_r;
logic din_ready_5_25;
logic din_almost_full_5_25;
logic [RID_WIDTH-1:0] hash_out_5_26;
logic hash_out_valid_filter_5_26;
rule_s_t din_5_26;
rule_s_t din_5_26_r1;
rule_s_t din_5_26_r2;
logic din_valid_5_26;
logic din_valid_5_26_r1;
logic din_valid_5_26_r2;
logic [2:0] din_valid_5_26_r;
logic din_ready_5_26;
logic din_almost_full_5_26;
logic [RID_WIDTH-1:0] hash_out_5_27;
logic hash_out_valid_filter_5_27;
rule_s_t din_5_27;
rule_s_t din_5_27_r1;
rule_s_t din_5_27_r2;
logic din_valid_5_27;
logic din_valid_5_27_r1;
logic din_valid_5_27_r2;
logic [2:0] din_valid_5_27_r;
logic din_ready_5_27;
logic din_almost_full_5_27;
logic [RID_WIDTH-1:0] hash_out_5_28;
logic hash_out_valid_filter_5_28;
rule_s_t din_5_28;
rule_s_t din_5_28_r1;
rule_s_t din_5_28_r2;
logic din_valid_5_28;
logic din_valid_5_28_r1;
logic din_valid_5_28_r2;
logic [2:0] din_valid_5_28_r;
logic din_ready_5_28;
logic din_almost_full_5_28;
logic [RID_WIDTH-1:0] hash_out_5_29;
logic hash_out_valid_filter_5_29;
rule_s_t din_5_29;
rule_s_t din_5_29_r1;
rule_s_t din_5_29_r2;
logic din_valid_5_29;
logic din_valid_5_29_r1;
logic din_valid_5_29_r2;
logic [2:0] din_valid_5_29_r;
logic din_ready_5_29;
logic din_almost_full_5_29;
logic [RID_WIDTH-1:0] hash_out_5_30;
logic hash_out_valid_filter_5_30;
rule_s_t din_5_30;
rule_s_t din_5_30_r1;
rule_s_t din_5_30_r2;
logic din_valid_5_30;
logic din_valid_5_30_r1;
logic din_valid_5_30_r2;
logic [2:0] din_valid_5_30_r;
logic din_ready_5_30;
logic din_almost_full_5_30;
logic [RID_WIDTH-1:0] hash_out_5_31;
logic hash_out_valid_filter_5_31;
rule_s_t din_5_31;
rule_s_t din_5_31_r1;
rule_s_t din_5_31_r2;
logic din_valid_5_31;
logic din_valid_5_31_r1;
logic din_valid_5_31_r2;
logic [2:0] din_valid_5_31_r;
logic din_ready_5_31;
logic din_almost_full_5_31;
logic [RID_WIDTH-1:0] hash_out_6_0;
logic hash_out_valid_filter_6_0;
rule_s_t din_6_0;
rule_s_t din_6_0_r1;
rule_s_t din_6_0_r2;
logic din_valid_6_0;
logic din_valid_6_0_r1;
logic din_valid_6_0_r2;
logic [2:0] din_valid_6_0_r;
logic din_ready_6_0;
logic din_almost_full_6_0;
logic [RID_WIDTH-1:0] hash_out_6_1;
logic hash_out_valid_filter_6_1;
rule_s_t din_6_1;
rule_s_t din_6_1_r1;
rule_s_t din_6_1_r2;
logic din_valid_6_1;
logic din_valid_6_1_r1;
logic din_valid_6_1_r2;
logic [2:0] din_valid_6_1_r;
logic din_ready_6_1;
logic din_almost_full_6_1;
logic [RID_WIDTH-1:0] hash_out_6_2;
logic hash_out_valid_filter_6_2;
rule_s_t din_6_2;
rule_s_t din_6_2_r1;
rule_s_t din_6_2_r2;
logic din_valid_6_2;
logic din_valid_6_2_r1;
logic din_valid_6_2_r2;
logic [2:0] din_valid_6_2_r;
logic din_ready_6_2;
logic din_almost_full_6_2;
logic [RID_WIDTH-1:0] hash_out_6_3;
logic hash_out_valid_filter_6_3;
rule_s_t din_6_3;
rule_s_t din_6_3_r1;
rule_s_t din_6_3_r2;
logic din_valid_6_3;
logic din_valid_6_3_r1;
logic din_valid_6_3_r2;
logic [2:0] din_valid_6_3_r;
logic din_ready_6_3;
logic din_almost_full_6_3;
logic [RID_WIDTH-1:0] hash_out_6_4;
logic hash_out_valid_filter_6_4;
rule_s_t din_6_4;
rule_s_t din_6_4_r1;
rule_s_t din_6_4_r2;
logic din_valid_6_4;
logic din_valid_6_4_r1;
logic din_valid_6_4_r2;
logic [2:0] din_valid_6_4_r;
logic din_ready_6_4;
logic din_almost_full_6_4;
logic [RID_WIDTH-1:0] hash_out_6_5;
logic hash_out_valid_filter_6_5;
rule_s_t din_6_5;
rule_s_t din_6_5_r1;
rule_s_t din_6_5_r2;
logic din_valid_6_5;
logic din_valid_6_5_r1;
logic din_valid_6_5_r2;
logic [2:0] din_valid_6_5_r;
logic din_ready_6_5;
logic din_almost_full_6_5;
logic [RID_WIDTH-1:0] hash_out_6_6;
logic hash_out_valid_filter_6_6;
rule_s_t din_6_6;
rule_s_t din_6_6_r1;
rule_s_t din_6_6_r2;
logic din_valid_6_6;
logic din_valid_6_6_r1;
logic din_valid_6_6_r2;
logic [2:0] din_valid_6_6_r;
logic din_ready_6_6;
logic din_almost_full_6_6;
logic [RID_WIDTH-1:0] hash_out_6_7;
logic hash_out_valid_filter_6_7;
rule_s_t din_6_7;
rule_s_t din_6_7_r1;
rule_s_t din_6_7_r2;
logic din_valid_6_7;
logic din_valid_6_7_r1;
logic din_valid_6_7_r2;
logic [2:0] din_valid_6_7_r;
logic din_ready_6_7;
logic din_almost_full_6_7;
logic [RID_WIDTH-1:0] hash_out_6_8;
logic hash_out_valid_filter_6_8;
rule_s_t din_6_8;
rule_s_t din_6_8_r1;
rule_s_t din_6_8_r2;
logic din_valid_6_8;
logic din_valid_6_8_r1;
logic din_valid_6_8_r2;
logic [2:0] din_valid_6_8_r;
logic din_ready_6_8;
logic din_almost_full_6_8;
logic [RID_WIDTH-1:0] hash_out_6_9;
logic hash_out_valid_filter_6_9;
rule_s_t din_6_9;
rule_s_t din_6_9_r1;
rule_s_t din_6_9_r2;
logic din_valid_6_9;
logic din_valid_6_9_r1;
logic din_valid_6_9_r2;
logic [2:0] din_valid_6_9_r;
logic din_ready_6_9;
logic din_almost_full_6_9;
logic [RID_WIDTH-1:0] hash_out_6_10;
logic hash_out_valid_filter_6_10;
rule_s_t din_6_10;
rule_s_t din_6_10_r1;
rule_s_t din_6_10_r2;
logic din_valid_6_10;
logic din_valid_6_10_r1;
logic din_valid_6_10_r2;
logic [2:0] din_valid_6_10_r;
logic din_ready_6_10;
logic din_almost_full_6_10;
logic [RID_WIDTH-1:0] hash_out_6_11;
logic hash_out_valid_filter_6_11;
rule_s_t din_6_11;
rule_s_t din_6_11_r1;
rule_s_t din_6_11_r2;
logic din_valid_6_11;
logic din_valid_6_11_r1;
logic din_valid_6_11_r2;
logic [2:0] din_valid_6_11_r;
logic din_ready_6_11;
logic din_almost_full_6_11;
logic [RID_WIDTH-1:0] hash_out_6_12;
logic hash_out_valid_filter_6_12;
rule_s_t din_6_12;
rule_s_t din_6_12_r1;
rule_s_t din_6_12_r2;
logic din_valid_6_12;
logic din_valid_6_12_r1;
logic din_valid_6_12_r2;
logic [2:0] din_valid_6_12_r;
logic din_ready_6_12;
logic din_almost_full_6_12;
logic [RID_WIDTH-1:0] hash_out_6_13;
logic hash_out_valid_filter_6_13;
rule_s_t din_6_13;
rule_s_t din_6_13_r1;
rule_s_t din_6_13_r2;
logic din_valid_6_13;
logic din_valid_6_13_r1;
logic din_valid_6_13_r2;
logic [2:0] din_valid_6_13_r;
logic din_ready_6_13;
logic din_almost_full_6_13;
logic [RID_WIDTH-1:0] hash_out_6_14;
logic hash_out_valid_filter_6_14;
rule_s_t din_6_14;
rule_s_t din_6_14_r1;
rule_s_t din_6_14_r2;
logic din_valid_6_14;
logic din_valid_6_14_r1;
logic din_valid_6_14_r2;
logic [2:0] din_valid_6_14_r;
logic din_ready_6_14;
logic din_almost_full_6_14;
logic [RID_WIDTH-1:0] hash_out_6_15;
logic hash_out_valid_filter_6_15;
rule_s_t din_6_15;
rule_s_t din_6_15_r1;
rule_s_t din_6_15_r2;
logic din_valid_6_15;
logic din_valid_6_15_r1;
logic din_valid_6_15_r2;
logic [2:0] din_valid_6_15_r;
logic din_ready_6_15;
logic din_almost_full_6_15;
logic [RID_WIDTH-1:0] hash_out_6_16;
logic hash_out_valid_filter_6_16;
rule_s_t din_6_16;
rule_s_t din_6_16_r1;
rule_s_t din_6_16_r2;
logic din_valid_6_16;
logic din_valid_6_16_r1;
logic din_valid_6_16_r2;
logic [2:0] din_valid_6_16_r;
logic din_ready_6_16;
logic din_almost_full_6_16;
logic [RID_WIDTH-1:0] hash_out_6_17;
logic hash_out_valid_filter_6_17;
rule_s_t din_6_17;
rule_s_t din_6_17_r1;
rule_s_t din_6_17_r2;
logic din_valid_6_17;
logic din_valid_6_17_r1;
logic din_valid_6_17_r2;
logic [2:0] din_valid_6_17_r;
logic din_ready_6_17;
logic din_almost_full_6_17;
logic [RID_WIDTH-1:0] hash_out_6_18;
logic hash_out_valid_filter_6_18;
rule_s_t din_6_18;
rule_s_t din_6_18_r1;
rule_s_t din_6_18_r2;
logic din_valid_6_18;
logic din_valid_6_18_r1;
logic din_valid_6_18_r2;
logic [2:0] din_valid_6_18_r;
logic din_ready_6_18;
logic din_almost_full_6_18;
logic [RID_WIDTH-1:0] hash_out_6_19;
logic hash_out_valid_filter_6_19;
rule_s_t din_6_19;
rule_s_t din_6_19_r1;
rule_s_t din_6_19_r2;
logic din_valid_6_19;
logic din_valid_6_19_r1;
logic din_valid_6_19_r2;
logic [2:0] din_valid_6_19_r;
logic din_ready_6_19;
logic din_almost_full_6_19;
logic [RID_WIDTH-1:0] hash_out_6_20;
logic hash_out_valid_filter_6_20;
rule_s_t din_6_20;
rule_s_t din_6_20_r1;
rule_s_t din_6_20_r2;
logic din_valid_6_20;
logic din_valid_6_20_r1;
logic din_valid_6_20_r2;
logic [2:0] din_valid_6_20_r;
logic din_ready_6_20;
logic din_almost_full_6_20;
logic [RID_WIDTH-1:0] hash_out_6_21;
logic hash_out_valid_filter_6_21;
rule_s_t din_6_21;
rule_s_t din_6_21_r1;
rule_s_t din_6_21_r2;
logic din_valid_6_21;
logic din_valid_6_21_r1;
logic din_valid_6_21_r2;
logic [2:0] din_valid_6_21_r;
logic din_ready_6_21;
logic din_almost_full_6_21;
logic [RID_WIDTH-1:0] hash_out_6_22;
logic hash_out_valid_filter_6_22;
rule_s_t din_6_22;
rule_s_t din_6_22_r1;
rule_s_t din_6_22_r2;
logic din_valid_6_22;
logic din_valid_6_22_r1;
logic din_valid_6_22_r2;
logic [2:0] din_valid_6_22_r;
logic din_ready_6_22;
logic din_almost_full_6_22;
logic [RID_WIDTH-1:0] hash_out_6_23;
logic hash_out_valid_filter_6_23;
rule_s_t din_6_23;
rule_s_t din_6_23_r1;
rule_s_t din_6_23_r2;
logic din_valid_6_23;
logic din_valid_6_23_r1;
logic din_valid_6_23_r2;
logic [2:0] din_valid_6_23_r;
logic din_ready_6_23;
logic din_almost_full_6_23;
logic [RID_WIDTH-1:0] hash_out_6_24;
logic hash_out_valid_filter_6_24;
rule_s_t din_6_24;
rule_s_t din_6_24_r1;
rule_s_t din_6_24_r2;
logic din_valid_6_24;
logic din_valid_6_24_r1;
logic din_valid_6_24_r2;
logic [2:0] din_valid_6_24_r;
logic din_ready_6_24;
logic din_almost_full_6_24;
logic [RID_WIDTH-1:0] hash_out_6_25;
logic hash_out_valid_filter_6_25;
rule_s_t din_6_25;
rule_s_t din_6_25_r1;
rule_s_t din_6_25_r2;
logic din_valid_6_25;
logic din_valid_6_25_r1;
logic din_valid_6_25_r2;
logic [2:0] din_valid_6_25_r;
logic din_ready_6_25;
logic din_almost_full_6_25;
logic [RID_WIDTH-1:0] hash_out_6_26;
logic hash_out_valid_filter_6_26;
rule_s_t din_6_26;
rule_s_t din_6_26_r1;
rule_s_t din_6_26_r2;
logic din_valid_6_26;
logic din_valid_6_26_r1;
logic din_valid_6_26_r2;
logic [2:0] din_valid_6_26_r;
logic din_ready_6_26;
logic din_almost_full_6_26;
logic [RID_WIDTH-1:0] hash_out_6_27;
logic hash_out_valid_filter_6_27;
rule_s_t din_6_27;
rule_s_t din_6_27_r1;
rule_s_t din_6_27_r2;
logic din_valid_6_27;
logic din_valid_6_27_r1;
logic din_valid_6_27_r2;
logic [2:0] din_valid_6_27_r;
logic din_ready_6_27;
logic din_almost_full_6_27;
logic [RID_WIDTH-1:0] hash_out_6_28;
logic hash_out_valid_filter_6_28;
rule_s_t din_6_28;
rule_s_t din_6_28_r1;
rule_s_t din_6_28_r2;
logic din_valid_6_28;
logic din_valid_6_28_r1;
logic din_valid_6_28_r2;
logic [2:0] din_valid_6_28_r;
logic din_ready_6_28;
logic din_almost_full_6_28;
logic [RID_WIDTH-1:0] hash_out_6_29;
logic hash_out_valid_filter_6_29;
rule_s_t din_6_29;
rule_s_t din_6_29_r1;
rule_s_t din_6_29_r2;
logic din_valid_6_29;
logic din_valid_6_29_r1;
logic din_valid_6_29_r2;
logic [2:0] din_valid_6_29_r;
logic din_ready_6_29;
logic din_almost_full_6_29;
logic [RID_WIDTH-1:0] hash_out_6_30;
logic hash_out_valid_filter_6_30;
rule_s_t din_6_30;
rule_s_t din_6_30_r1;
rule_s_t din_6_30_r2;
logic din_valid_6_30;
logic din_valid_6_30_r1;
logic din_valid_6_30_r2;
logic [2:0] din_valid_6_30_r;
logic din_ready_6_30;
logic din_almost_full_6_30;
logic [RID_WIDTH-1:0] hash_out_6_31;
logic hash_out_valid_filter_6_31;
rule_s_t din_6_31;
rule_s_t din_6_31_r1;
rule_s_t din_6_31_r2;
logic din_valid_6_31;
logic din_valid_6_31_r1;
logic din_valid_6_31_r2;
logic [2:0] din_valid_6_31_r;
logic din_ready_6_31;
logic din_almost_full_6_31;
logic [RID_WIDTH-1:0] hash_out_7_0;
logic hash_out_valid_filter_7_0;
rule_s_t din_7_0;
rule_s_t din_7_0_r1;
rule_s_t din_7_0_r2;
logic din_valid_7_0;
logic din_valid_7_0_r1;
logic din_valid_7_0_r2;
logic [2:0] din_valid_7_0_r;
logic din_ready_7_0;
logic din_almost_full_7_0;
logic [RID_WIDTH-1:0] hash_out_7_1;
logic hash_out_valid_filter_7_1;
rule_s_t din_7_1;
rule_s_t din_7_1_r1;
rule_s_t din_7_1_r2;
logic din_valid_7_1;
logic din_valid_7_1_r1;
logic din_valid_7_1_r2;
logic [2:0] din_valid_7_1_r;
logic din_ready_7_1;
logic din_almost_full_7_1;
logic [RID_WIDTH-1:0] hash_out_7_2;
logic hash_out_valid_filter_7_2;
rule_s_t din_7_2;
rule_s_t din_7_2_r1;
rule_s_t din_7_2_r2;
logic din_valid_7_2;
logic din_valid_7_2_r1;
logic din_valid_7_2_r2;
logic [2:0] din_valid_7_2_r;
logic din_ready_7_2;
logic din_almost_full_7_2;
logic [RID_WIDTH-1:0] hash_out_7_3;
logic hash_out_valid_filter_7_3;
rule_s_t din_7_3;
rule_s_t din_7_3_r1;
rule_s_t din_7_3_r2;
logic din_valid_7_3;
logic din_valid_7_3_r1;
logic din_valid_7_3_r2;
logic [2:0] din_valid_7_3_r;
logic din_ready_7_3;
logic din_almost_full_7_3;
logic [RID_WIDTH-1:0] hash_out_7_4;
logic hash_out_valid_filter_7_4;
rule_s_t din_7_4;
rule_s_t din_7_4_r1;
rule_s_t din_7_4_r2;
logic din_valid_7_4;
logic din_valid_7_4_r1;
logic din_valid_7_4_r2;
logic [2:0] din_valid_7_4_r;
logic din_ready_7_4;
logic din_almost_full_7_4;
logic [RID_WIDTH-1:0] hash_out_7_5;
logic hash_out_valid_filter_7_5;
rule_s_t din_7_5;
rule_s_t din_7_5_r1;
rule_s_t din_7_5_r2;
logic din_valid_7_5;
logic din_valid_7_5_r1;
logic din_valid_7_5_r2;
logic [2:0] din_valid_7_5_r;
logic din_ready_7_5;
logic din_almost_full_7_5;
logic [RID_WIDTH-1:0] hash_out_7_6;
logic hash_out_valid_filter_7_6;
rule_s_t din_7_6;
rule_s_t din_7_6_r1;
rule_s_t din_7_6_r2;
logic din_valid_7_6;
logic din_valid_7_6_r1;
logic din_valid_7_6_r2;
logic [2:0] din_valid_7_6_r;
logic din_ready_7_6;
logic din_almost_full_7_6;
logic [RID_WIDTH-1:0] hash_out_7_7;
logic hash_out_valid_filter_7_7;
rule_s_t din_7_7;
rule_s_t din_7_7_r1;
rule_s_t din_7_7_r2;
logic din_valid_7_7;
logic din_valid_7_7_r1;
logic din_valid_7_7_r2;
logic [2:0] din_valid_7_7_r;
logic din_ready_7_7;
logic din_almost_full_7_7;
logic [RID_WIDTH-1:0] hash_out_7_8;
logic hash_out_valid_filter_7_8;
rule_s_t din_7_8;
rule_s_t din_7_8_r1;
rule_s_t din_7_8_r2;
logic din_valid_7_8;
logic din_valid_7_8_r1;
logic din_valid_7_8_r2;
logic [2:0] din_valid_7_8_r;
logic din_ready_7_8;
logic din_almost_full_7_8;
logic [RID_WIDTH-1:0] hash_out_7_9;
logic hash_out_valid_filter_7_9;
rule_s_t din_7_9;
rule_s_t din_7_9_r1;
rule_s_t din_7_9_r2;
logic din_valid_7_9;
logic din_valid_7_9_r1;
logic din_valid_7_9_r2;
logic [2:0] din_valid_7_9_r;
logic din_ready_7_9;
logic din_almost_full_7_9;
logic [RID_WIDTH-1:0] hash_out_7_10;
logic hash_out_valid_filter_7_10;
rule_s_t din_7_10;
rule_s_t din_7_10_r1;
rule_s_t din_7_10_r2;
logic din_valid_7_10;
logic din_valid_7_10_r1;
logic din_valid_7_10_r2;
logic [2:0] din_valid_7_10_r;
logic din_ready_7_10;
logic din_almost_full_7_10;
logic [RID_WIDTH-1:0] hash_out_7_11;
logic hash_out_valid_filter_7_11;
rule_s_t din_7_11;
rule_s_t din_7_11_r1;
rule_s_t din_7_11_r2;
logic din_valid_7_11;
logic din_valid_7_11_r1;
logic din_valid_7_11_r2;
logic [2:0] din_valid_7_11_r;
logic din_ready_7_11;
logic din_almost_full_7_11;
logic [RID_WIDTH-1:0] hash_out_7_12;
logic hash_out_valid_filter_7_12;
rule_s_t din_7_12;
rule_s_t din_7_12_r1;
rule_s_t din_7_12_r2;
logic din_valid_7_12;
logic din_valid_7_12_r1;
logic din_valid_7_12_r2;
logic [2:0] din_valid_7_12_r;
logic din_ready_7_12;
logic din_almost_full_7_12;
logic [RID_WIDTH-1:0] hash_out_7_13;
logic hash_out_valid_filter_7_13;
rule_s_t din_7_13;
rule_s_t din_7_13_r1;
rule_s_t din_7_13_r2;
logic din_valid_7_13;
logic din_valid_7_13_r1;
logic din_valid_7_13_r2;
logic [2:0] din_valid_7_13_r;
logic din_ready_7_13;
logic din_almost_full_7_13;
logic [RID_WIDTH-1:0] hash_out_7_14;
logic hash_out_valid_filter_7_14;
rule_s_t din_7_14;
rule_s_t din_7_14_r1;
rule_s_t din_7_14_r2;
logic din_valid_7_14;
logic din_valid_7_14_r1;
logic din_valid_7_14_r2;
logic [2:0] din_valid_7_14_r;
logic din_ready_7_14;
logic din_almost_full_7_14;
logic [RID_WIDTH-1:0] hash_out_7_15;
logic hash_out_valid_filter_7_15;
rule_s_t din_7_15;
rule_s_t din_7_15_r1;
rule_s_t din_7_15_r2;
logic din_valid_7_15;
logic din_valid_7_15_r1;
logic din_valid_7_15_r2;
logic [2:0] din_valid_7_15_r;
logic din_ready_7_15;
logic din_almost_full_7_15;
logic [RID_WIDTH-1:0] hash_out_7_16;
logic hash_out_valid_filter_7_16;
rule_s_t din_7_16;
rule_s_t din_7_16_r1;
rule_s_t din_7_16_r2;
logic din_valid_7_16;
logic din_valid_7_16_r1;
logic din_valid_7_16_r2;
logic [2:0] din_valid_7_16_r;
logic din_ready_7_16;
logic din_almost_full_7_16;
logic [RID_WIDTH-1:0] hash_out_7_17;
logic hash_out_valid_filter_7_17;
rule_s_t din_7_17;
rule_s_t din_7_17_r1;
rule_s_t din_7_17_r2;
logic din_valid_7_17;
logic din_valid_7_17_r1;
logic din_valid_7_17_r2;
logic [2:0] din_valid_7_17_r;
logic din_ready_7_17;
logic din_almost_full_7_17;
logic [RID_WIDTH-1:0] hash_out_7_18;
logic hash_out_valid_filter_7_18;
rule_s_t din_7_18;
rule_s_t din_7_18_r1;
rule_s_t din_7_18_r2;
logic din_valid_7_18;
logic din_valid_7_18_r1;
logic din_valid_7_18_r2;
logic [2:0] din_valid_7_18_r;
logic din_ready_7_18;
logic din_almost_full_7_18;
logic [RID_WIDTH-1:0] hash_out_7_19;
logic hash_out_valid_filter_7_19;
rule_s_t din_7_19;
rule_s_t din_7_19_r1;
rule_s_t din_7_19_r2;
logic din_valid_7_19;
logic din_valid_7_19_r1;
logic din_valid_7_19_r2;
logic [2:0] din_valid_7_19_r;
logic din_ready_7_19;
logic din_almost_full_7_19;
logic [RID_WIDTH-1:0] hash_out_7_20;
logic hash_out_valid_filter_7_20;
rule_s_t din_7_20;
rule_s_t din_7_20_r1;
rule_s_t din_7_20_r2;
logic din_valid_7_20;
logic din_valid_7_20_r1;
logic din_valid_7_20_r2;
logic [2:0] din_valid_7_20_r;
logic din_ready_7_20;
logic din_almost_full_7_20;
logic [RID_WIDTH-1:0] hash_out_7_21;
logic hash_out_valid_filter_7_21;
rule_s_t din_7_21;
rule_s_t din_7_21_r1;
rule_s_t din_7_21_r2;
logic din_valid_7_21;
logic din_valid_7_21_r1;
logic din_valid_7_21_r2;
logic [2:0] din_valid_7_21_r;
logic din_ready_7_21;
logic din_almost_full_7_21;
logic [RID_WIDTH-1:0] hash_out_7_22;
logic hash_out_valid_filter_7_22;
rule_s_t din_7_22;
rule_s_t din_7_22_r1;
rule_s_t din_7_22_r2;
logic din_valid_7_22;
logic din_valid_7_22_r1;
logic din_valid_7_22_r2;
logic [2:0] din_valid_7_22_r;
logic din_ready_7_22;
logic din_almost_full_7_22;
logic [RID_WIDTH-1:0] hash_out_7_23;
logic hash_out_valid_filter_7_23;
rule_s_t din_7_23;
rule_s_t din_7_23_r1;
rule_s_t din_7_23_r2;
logic din_valid_7_23;
logic din_valid_7_23_r1;
logic din_valid_7_23_r2;
logic [2:0] din_valid_7_23_r;
logic din_ready_7_23;
logic din_almost_full_7_23;
logic [RID_WIDTH-1:0] hash_out_7_24;
logic hash_out_valid_filter_7_24;
rule_s_t din_7_24;
rule_s_t din_7_24_r1;
rule_s_t din_7_24_r2;
logic din_valid_7_24;
logic din_valid_7_24_r1;
logic din_valid_7_24_r2;
logic [2:0] din_valid_7_24_r;
logic din_ready_7_24;
logic din_almost_full_7_24;
logic [RID_WIDTH-1:0] hash_out_7_25;
logic hash_out_valid_filter_7_25;
rule_s_t din_7_25;
rule_s_t din_7_25_r1;
rule_s_t din_7_25_r2;
logic din_valid_7_25;
logic din_valid_7_25_r1;
logic din_valid_7_25_r2;
logic [2:0] din_valid_7_25_r;
logic din_ready_7_25;
logic din_almost_full_7_25;
logic [RID_WIDTH-1:0] hash_out_7_26;
logic hash_out_valid_filter_7_26;
rule_s_t din_7_26;
rule_s_t din_7_26_r1;
rule_s_t din_7_26_r2;
logic din_valid_7_26;
logic din_valid_7_26_r1;
logic din_valid_7_26_r2;
logic [2:0] din_valid_7_26_r;
logic din_ready_7_26;
logic din_almost_full_7_26;
logic [RID_WIDTH-1:0] hash_out_7_27;
logic hash_out_valid_filter_7_27;
rule_s_t din_7_27;
rule_s_t din_7_27_r1;
rule_s_t din_7_27_r2;
logic din_valid_7_27;
logic din_valid_7_27_r1;
logic din_valid_7_27_r2;
logic [2:0] din_valid_7_27_r;
logic din_ready_7_27;
logic din_almost_full_7_27;
logic [RID_WIDTH-1:0] hash_out_7_28;
logic hash_out_valid_filter_7_28;
rule_s_t din_7_28;
rule_s_t din_7_28_r1;
rule_s_t din_7_28_r2;
logic din_valid_7_28;
logic din_valid_7_28_r1;
logic din_valid_7_28_r2;
logic [2:0] din_valid_7_28_r;
logic din_ready_7_28;
logic din_almost_full_7_28;
logic [RID_WIDTH-1:0] hash_out_7_29;
logic hash_out_valid_filter_7_29;
rule_s_t din_7_29;
rule_s_t din_7_29_r1;
rule_s_t din_7_29_r2;
logic din_valid_7_29;
logic din_valid_7_29_r1;
logic din_valid_7_29_r2;
logic [2:0] din_valid_7_29_r;
logic din_ready_7_29;
logic din_almost_full_7_29;
logic [RID_WIDTH-1:0] hash_out_7_30;
logic hash_out_valid_filter_7_30;
rule_s_t din_7_30;
rule_s_t din_7_30_r1;
rule_s_t din_7_30_r2;
logic din_valid_7_30;
logic din_valid_7_30_r1;
logic din_valid_7_30_r2;
logic [2:0] din_valid_7_30_r;
logic din_ready_7_30;
logic din_almost_full_7_30;
logic [RID_WIDTH-1:0] hash_out_7_31;
logic hash_out_valid_filter_7_31;
rule_s_t din_7_31;
rule_s_t din_7_31_r1;
rule_s_t din_7_31_r2;
logic din_valid_7_31;
logic din_valid_7_31_r1;
logic din_valid_7_31_r2;
logic [2:0] din_valid_7_31_r;
logic din_ready_7_31;
logic din_almost_full_7_31;

logic out_new_pkt;

logic [255:0] in_convt;
logic gap;

//status 
logic [7:0] status_addr_r;
logic [STAT_AWIDTH-1:0]  status_addr_sel_r;
logic status_write_r;
logic status_read_r;
logic [31:0] status_writedata_r;
logic [31:0] status_readdata_sm;
logic status_readdata_valid_sm;
logic [31:0] status_readdata_back;
logic status_readdata_valid_back;
logic [31:0] test_valid_cnt = 0;
logic [31:0] test_empty;
logic [31:0] test_din_0;
logic [31:0] test_din_r2_0;
logic [31:0] test_din_1;
logic [31:0] test_din_r2_1;
logic [31:0] test_din_2;
logic [31:0] test_din_r2_2;
logic [31:0] test_din_3;
logic [31:0] test_din_r2_3;
logic [31:0] test_din_4;
logic [31:0] test_din_r2_4;
logic [31:0] test_din_5;
logic [31:0] test_din_r2_5;
logic [31:0] test_din_6;
logic [31:0] test_din_r2_6;
logic [31:0] test_din_7;
logic [31:0] test_din_r2_7;

assign in_convt[7+0*8:0+0*8] = in_data[255-0*8:255-7-0*8];
assign in_convt[7+1*8:0+1*8] = in_data[255-1*8:255-7-1*8];
assign in_convt[7+2*8:0+2*8] = in_data[255-2*8:255-7-2*8];
assign in_convt[7+3*8:0+3*8] = in_data[255-3*8:255-7-3*8];
assign in_convt[7+4*8:0+4*8] = in_data[255-4*8:255-7-4*8];
assign in_convt[7+5*8:0+5*8] = in_data[255-5*8:255-7-5*8];
assign in_convt[7+6*8:0+6*8] = in_data[255-6*8:255-7-6*8];
assign in_convt[7+7*8:0+7*8] = in_data[255-7*8:255-7-7*8];
assign in_convt[7+8*8:0+8*8] = in_data[255-8*8:255-7-8*8];
assign in_convt[7+9*8:0+9*8] = in_data[255-9*8:255-7-9*8];
assign in_convt[7+10*8:0+10*8] = in_data[255-10*8:255-7-10*8];
assign in_convt[7+11*8:0+11*8] = in_data[255-11*8:255-7-11*8];
assign in_convt[7+12*8:0+12*8] = in_data[255-12*8:255-7-12*8];
assign in_convt[7+13*8:0+13*8] = in_data[255-13*8:255-7-13*8];
assign in_convt[7+14*8:0+14*8] = in_data[255-14*8:255-7-14*8];
assign in_convt[7+15*8:0+15*8] = in_data[255-15*8:255-7-15*8];
assign in_convt[7+16*8:0+16*8] = in_data[255-16*8:255-7-16*8];
assign in_convt[7+17*8:0+17*8] = in_data[255-17*8:255-7-17*8];
assign in_convt[7+18*8:0+18*8] = in_data[255-18*8:255-7-18*8];
assign in_convt[7+19*8:0+19*8] = in_data[255-19*8:255-7-19*8];
assign in_convt[7+20*8:0+20*8] = in_data[255-20*8:255-7-20*8];
assign in_convt[7+21*8:0+21*8] = in_data[255-21*8:255-7-21*8];
assign in_convt[7+22*8:0+22*8] = in_data[255-22*8:255-7-22*8];
assign in_convt[7+23*8:0+23*8] = in_data[255-23*8:255-7-23*8];
assign in_convt[7+24*8:0+24*8] = in_data[255-24*8:255-7-24*8];
assign in_convt[7+25*8:0+25*8] = in_data[255-25*8:255-7-25*8];
assign in_convt[7+26*8:0+26*8] = in_data[255-26*8:255-7-26*8];
assign in_convt[7+27*8:0+27*8] = in_data[255-27*8:255-7-27*8];
assign in_convt[7+28*8:0+28*8] = in_data[255-28*8:255-7-28*8];
assign in_convt[7+29*8:0+29*8] = in_data[255-29*8:255-7-29*8];
assign in_convt[7+30*8:0+30*8] = in_data[255-30*8:255-7-30*8];
assign in_convt[7+31*8:0+31*8] = in_data[255-31*8:255-7-31*8];

always @ (posedge clk) begin
    //in_ready <=   !din_almost_full_0_0 &  !din_almost_full_0_1 &  !din_almost_full_0_2 &  !din_almost_full_0_3 &  !din_almost_full_0_4 &  !din_almost_full_0_5 &  !din_almost_full_0_6 &  !din_almost_full_0_7 &  !din_almost_full_0_8 &  !din_almost_full_0_9 &  !din_almost_full_0_10 &  !din_almost_full_0_11 &  !din_almost_full_0_12 &  !din_almost_full_0_13 &  !din_almost_full_0_14 &  !din_almost_full_0_15 &  !din_almost_full_0_16 &  !din_almost_full_0_17 &  !din_almost_full_0_18 &  !din_almost_full_0_19 &  !din_almost_full_0_20 &  !din_almost_full_0_21 &  !din_almost_full_0_22 &  !din_almost_full_0_23 &  !din_almost_full_0_24 &  !din_almost_full_0_25 &  !din_almost_full_0_26 &  !din_almost_full_0_27 &  !din_almost_full_0_28 &  !din_almost_full_0_29 &  !din_almost_full_0_30 &  !din_almost_full_0_31 &    !din_almost_full_1_0 &  !din_almost_full_1_1 &  !din_almost_full_1_2 &  !din_almost_full_1_3 &  !din_almost_full_1_4 &  !din_almost_full_1_5 &  !din_almost_full_1_6 &  !din_almost_full_1_7 &  !din_almost_full_1_8 &  !din_almost_full_1_9 &  !din_almost_full_1_10 &  !din_almost_full_1_11 &  !din_almost_full_1_12 &  !din_almost_full_1_13 &  !din_almost_full_1_14 &  !din_almost_full_1_15 &  !din_almost_full_1_16 &  !din_almost_full_1_17 &  !din_almost_full_1_18 &  !din_almost_full_1_19 &  !din_almost_full_1_20 &  !din_almost_full_1_21 &  !din_almost_full_1_22 &  !din_almost_full_1_23 &  !din_almost_full_1_24 &  !din_almost_full_1_25 &  !din_almost_full_1_26 &  !din_almost_full_1_27 &  !din_almost_full_1_28 &  !din_almost_full_1_29 &  !din_almost_full_1_30 &  !din_almost_full_1_31 &    !din_almost_full_2_0 &  !din_almost_full_2_1 &  !din_almost_full_2_2 &  !din_almost_full_2_3 &  !din_almost_full_2_4 &  !din_almost_full_2_5 &  !din_almost_full_2_6 &  !din_almost_full_2_7 &  !din_almost_full_2_8 &  !din_almost_full_2_9 &  !din_almost_full_2_10 &  !din_almost_full_2_11 &  !din_almost_full_2_12 &  !din_almost_full_2_13 &  !din_almost_full_2_14 &  !din_almost_full_2_15 &  !din_almost_full_2_16 &  !din_almost_full_2_17 &  !din_almost_full_2_18 &  !din_almost_full_2_19 &  !din_almost_full_2_20 &  !din_almost_full_2_21 &  !din_almost_full_2_22 &  !din_almost_full_2_23 &  !din_almost_full_2_24 &  !din_almost_full_2_25 &  !din_almost_full_2_26 &  !din_almost_full_2_27 &  !din_almost_full_2_28 &  !din_almost_full_2_29 &  !din_almost_full_2_30 &  !din_almost_full_2_31 &    !din_almost_full_3_0 &  !din_almost_full_3_1 &  !din_almost_full_3_2 &  !din_almost_full_3_3 &  !din_almost_full_3_4 &  !din_almost_full_3_5 &  !din_almost_full_3_6 &  !din_almost_full_3_7 &  !din_almost_full_3_8 &  !din_almost_full_3_9 &  !din_almost_full_3_10 &  !din_almost_full_3_11 &  !din_almost_full_3_12 &  !din_almost_full_3_13 &  !din_almost_full_3_14 &  !din_almost_full_3_15 &  !din_almost_full_3_16 &  !din_almost_full_3_17 &  !din_almost_full_3_18 &  !din_almost_full_3_19 &  !din_almost_full_3_20 &  !din_almost_full_3_21 &  !din_almost_full_3_22 &  !din_almost_full_3_23 &  !din_almost_full_3_24 &  !din_almost_full_3_25 &  !din_almost_full_3_26 &  !din_almost_full_3_27 &  !din_almost_full_3_28 &  !din_almost_full_3_29 &  !din_almost_full_3_30 &  !din_almost_full_3_31 &    !din_almost_full_4_0 &  !din_almost_full_4_1 &  !din_almost_full_4_2 &  !din_almost_full_4_3 &  !din_almost_full_4_4 &  !din_almost_full_4_5 &  !din_almost_full_4_6 &  !din_almost_full_4_7 &  !din_almost_full_4_8 &  !din_almost_full_4_9 &  !din_almost_full_4_10 &  !din_almost_full_4_11 &  !din_almost_full_4_12 &  !din_almost_full_4_13 &  !din_almost_full_4_14 &  !din_almost_full_4_15 &  !din_almost_full_4_16 &  !din_almost_full_4_17 &  !din_almost_full_4_18 &  !din_almost_full_4_19 &  !din_almost_full_4_20 &  !din_almost_full_4_21 &  !din_almost_full_4_22 &  !din_almost_full_4_23 &  !din_almost_full_4_24 &  !din_almost_full_4_25 &  !din_almost_full_4_26 &  !din_almost_full_4_27 &  !din_almost_full_4_28 &  !din_almost_full_4_29 &  !din_almost_full_4_30 &  !din_almost_full_4_31 &    !din_almost_full_5_0 &  !din_almost_full_5_1 &  !din_almost_full_5_2 &  !din_almost_full_5_3 &  !din_almost_full_5_4 &  !din_almost_full_5_5 &  !din_almost_full_5_6 &  !din_almost_full_5_7 &  !din_almost_full_5_8 &  !din_almost_full_5_9 &  !din_almost_full_5_10 &  !din_almost_full_5_11 &  !din_almost_full_5_12 &  !din_almost_full_5_13 &  !din_almost_full_5_14 &  !din_almost_full_5_15 &  !din_almost_full_5_16 &  !din_almost_full_5_17 &  !din_almost_full_5_18 &  !din_almost_full_5_19 &  !din_almost_full_5_20 &  !din_almost_full_5_21 &  !din_almost_full_5_22 &  !din_almost_full_5_23 &  !din_almost_full_5_24 &  !din_almost_full_5_25 &  !din_almost_full_5_26 &  !din_almost_full_5_27 &  !din_almost_full_5_28 &  !din_almost_full_5_29 &  !din_almost_full_5_30 &  !din_almost_full_5_31 &    !din_almost_full_6_0 &  !din_almost_full_6_1 &  !din_almost_full_6_2 &  !din_almost_full_6_3 &  !din_almost_full_6_4 &  !din_almost_full_6_5 &  !din_almost_full_6_6 &  !din_almost_full_6_7 &  !din_almost_full_6_8 &  !din_almost_full_6_9 &  !din_almost_full_6_10 &  !din_almost_full_6_11 &  !din_almost_full_6_12 &  !din_almost_full_6_13 &  !din_almost_full_6_14 &  !din_almost_full_6_15 &  !din_almost_full_6_16 &  !din_almost_full_6_17 &  !din_almost_full_6_18 &  !din_almost_full_6_19 &  !din_almost_full_6_20 &  !din_almost_full_6_21 &  !din_almost_full_6_22 &  !din_almost_full_6_23 &  !din_almost_full_6_24 &  !din_almost_full_6_25 &  !din_almost_full_6_26 &  !din_almost_full_6_27 &  !din_almost_full_6_28 &  !din_almost_full_6_29 &  !din_almost_full_6_30 &  !din_almost_full_6_31 &    !din_almost_full_7_0 &  !din_almost_full_7_1 &  !din_almost_full_7_2 &  !din_almost_full_7_3 &  !din_almost_full_7_4 &  !din_almost_full_7_5 &  !din_almost_full_7_6 &  !din_almost_full_7_7 &  !din_almost_full_7_8 &  !din_almost_full_7_9 &  !din_almost_full_7_10 &  !din_almost_full_7_11 &  !din_almost_full_7_12 &  !din_almost_full_7_13 &  !din_almost_full_7_14 &  !din_almost_full_7_15 &  !din_almost_full_7_16 &  !din_almost_full_7_17 &  !din_almost_full_7_18 &  !din_almost_full_7_19 &  !din_almost_full_7_20 &  !din_almost_full_7_21 &  !din_almost_full_7_22 &  !din_almost_full_7_23 &  !din_almost_full_7_24 &  !din_almost_full_7_25 &  !din_almost_full_7_26 &  !din_almost_full_7_27 &  !din_almost_full_7_28 &  !din_almost_full_7_29 &  !din_almost_full_7_30 &  !din_almost_full_7_31 &   !gap;
    in_ready <=   !din_almost_full_0_0 &  !din_almost_full_0_1 &  !din_almost_full_0_2 &  !din_almost_full_0_3 &  !din_almost_full_0_4 &  !din_almost_full_0_5 &  !din_almost_full_0_6 &  !din_almost_full_0_7 &  !din_almost_full_0_8 &  !din_almost_full_0_9 &  !din_almost_full_0_10 &  !din_almost_full_0_11 &  !din_almost_full_0_12 &  !din_almost_full_0_13 &  !din_almost_full_0_14 &  !din_almost_full_0_15 &  !din_almost_full_0_16 &  !din_almost_full_0_17 &  !din_almost_full_0_18 &  !din_almost_full_0_19 &  !din_almost_full_0_20 &  !din_almost_full_0_21 &  !din_almost_full_0_22 &  !din_almost_full_0_23 &  !din_almost_full_0_24 &  !din_almost_full_0_25 &  !din_almost_full_0_26 &  !din_almost_full_0_27 &  !din_almost_full_0_28 &  !din_almost_full_0_29 &  !din_almost_full_0_30 &  !din_almost_full_0_31 &    !din_almost_full_1_0 &  !din_almost_full_1_1 &  !din_almost_full_1_2 &  !din_almost_full_1_3 &  !din_almost_full_1_4 &  !din_almost_full_1_5 &  !din_almost_full_1_6 &  !din_almost_full_1_7 &  !din_almost_full_1_8 &  !din_almost_full_1_9 &  !din_almost_full_1_10 &  !din_almost_full_1_11 &  !din_almost_full_1_12 &  !din_almost_full_1_13 &  !din_almost_full_1_14 &  !din_almost_full_1_15 &  !din_almost_full_1_16 &  !din_almost_full_1_17 &  !din_almost_full_1_18 &  !din_almost_full_1_19 &  !din_almost_full_1_20 &  !din_almost_full_1_21 &  !din_almost_full_1_22 &  !din_almost_full_1_23 &  !din_almost_full_1_24 &  !din_almost_full_1_25 &  !din_almost_full_1_26 &  !din_almost_full_1_27 &  !din_almost_full_1_28 &  !din_almost_full_1_29 &  !din_almost_full_1_30 &  !din_almost_full_1_31 &    !din_almost_full_2_0 &  !din_almost_full_2_1 &  !din_almost_full_2_2 &  !din_almost_full_2_3 &  !din_almost_full_2_4 &  !din_almost_full_2_5 &  !din_almost_full_2_6 &  !din_almost_full_2_7 &  !din_almost_full_2_8 &  !din_almost_full_2_9 &  !din_almost_full_2_10 &  !din_almost_full_2_11 &  !din_almost_full_2_12 &  !din_almost_full_2_13 &  !din_almost_full_2_14 &  !din_almost_full_2_15 &  !din_almost_full_2_16 &  !din_almost_full_2_17 &  !din_almost_full_2_18 &  !din_almost_full_2_19 &  !din_almost_full_2_20 &  !din_almost_full_2_21 &  !din_almost_full_2_22 &  !din_almost_full_2_23 &  !din_almost_full_2_24 &  !din_almost_full_2_25 &  !din_almost_full_2_26 &  !din_almost_full_2_27 &  !din_almost_full_2_28 &  !din_almost_full_2_29 &  !din_almost_full_2_30 &  !din_almost_full_2_31 &    !din_almost_full_3_0 &  !din_almost_full_3_1 &  !din_almost_full_3_2 &  !din_almost_full_3_3 &  !din_almost_full_3_4 &  !din_almost_full_3_5 &  !din_almost_full_3_6 &  !din_almost_full_3_7 &  !din_almost_full_3_8 &  !din_almost_full_3_9 &  !din_almost_full_3_10 &  !din_almost_full_3_11 &  !din_almost_full_3_12 &  !din_almost_full_3_13 &  !din_almost_full_3_14 &  !din_almost_full_3_15 &  !din_almost_full_3_16 &  !din_almost_full_3_17 &  !din_almost_full_3_18 &  !din_almost_full_3_19 &  !din_almost_full_3_20 &  !din_almost_full_3_21 &  !din_almost_full_3_22 &  !din_almost_full_3_23 &  !din_almost_full_3_24 &  !din_almost_full_3_25 &  !din_almost_full_3_26 &  !din_almost_full_3_27 &  !din_almost_full_3_28 &  !din_almost_full_3_29 &  !din_almost_full_3_30 &  !din_almost_full_3_31 &    !din_almost_full_4_0 &  !din_almost_full_4_1 &  !din_almost_full_4_2 &  !din_almost_full_4_3 &  !din_almost_full_4_4 &  !din_almost_full_4_5 &  !din_almost_full_4_6 &  !din_almost_full_4_7 &  !din_almost_full_4_8 &  !din_almost_full_4_9 &  !din_almost_full_4_10 &  !din_almost_full_4_11 &  !din_almost_full_4_12 &  !din_almost_full_4_13 &  !din_almost_full_4_14 &  !din_almost_full_4_15 &  !din_almost_full_4_16 &  !din_almost_full_4_17 &  !din_almost_full_4_18 &  !din_almost_full_4_19 &  !din_almost_full_4_20 &  !din_almost_full_4_21 &  !din_almost_full_4_22 &  !din_almost_full_4_23 &  !din_almost_full_4_24 &  !din_almost_full_4_25 &  !din_almost_full_4_26 &  !din_almost_full_4_27 &  !din_almost_full_4_28 &  !din_almost_full_4_29 &  !din_almost_full_4_30 &  !din_almost_full_4_31 &    !din_almost_full_5_0 &  !din_almost_full_5_1 &  !din_almost_full_5_2 &  !din_almost_full_5_3 &  !din_almost_full_5_4 &  !din_almost_full_5_5 &  !din_almost_full_5_6 &  !din_almost_full_5_7 &  !din_almost_full_5_8 &  !din_almost_full_5_9 &  !din_almost_full_5_10 &  !din_almost_full_5_11 &  !din_almost_full_5_12 &  !din_almost_full_5_13 &  !din_almost_full_5_14 &  !din_almost_full_5_15 &  !din_almost_full_5_16 &  !din_almost_full_5_17 &  !din_almost_full_5_18 &  !din_almost_full_5_19 &  !din_almost_full_5_20 &  !din_almost_full_5_21 &  !din_almost_full_5_22 &  !din_almost_full_5_23 &  !din_almost_full_5_24 &  !din_almost_full_5_25 &  !din_almost_full_5_26 &  !din_almost_full_5_27 &  !din_almost_full_5_28 &  !din_almost_full_5_29 &  !din_almost_full_5_30 &  !din_almost_full_5_31 &    !din_almost_full_6_0 &  !din_almost_full_6_1 &  !din_almost_full_6_2 &  !din_almost_full_6_3 &  !din_almost_full_6_4 &  !din_almost_full_6_5 &  !din_almost_full_6_6 &  !din_almost_full_6_7 &  !din_almost_full_6_8 &  !din_almost_full_6_9 &  !din_almost_full_6_10 &  !din_almost_full_6_11 &  !din_almost_full_6_12 &  !din_almost_full_6_13 &  !din_almost_full_6_14 &  !din_almost_full_6_15 &  !din_almost_full_6_16 &  !din_almost_full_6_17 &  !din_almost_full_6_18 &  !din_almost_full_6_19 &  !din_almost_full_6_20 &  !din_almost_full_6_21 &  !din_almost_full_6_22 &  !din_almost_full_6_23 &  !din_almost_full_6_24 &  !din_almost_full_6_25 &  !din_almost_full_6_26 &  !din_almost_full_6_27 &  !din_almost_full_6_28 &  !din_almost_full_6_29 &  !din_almost_full_6_30 &  !din_almost_full_6_31 &    !din_almost_full_7_0 &  !din_almost_full_7_1 &  !din_almost_full_7_2 &  !din_almost_full_7_3 &  !din_almost_full_7_4 &  !din_almost_full_7_5 &  !din_almost_full_7_6 &  !din_almost_full_7_7 &  !din_almost_full_7_8 &  !din_almost_full_7_9 &  !din_almost_full_7_10 &  !din_almost_full_7_11 &  !din_almost_full_7_12 &  !din_almost_full_7_13 &  !din_almost_full_7_14 &  !din_almost_full_7_15 &  !din_almost_full_7_16 &  !din_almost_full_7_17 &  !din_almost_full_7_18 &  !din_almost_full_7_19 &  !din_almost_full_7_20 &  !din_almost_full_7_21 &  !din_almost_full_7_22 &  !din_almost_full_7_23 &  !din_almost_full_7_24 &  !din_almost_full_7_25 &  !din_almost_full_7_26 &  !din_almost_full_7_27 &  !din_almost_full_7_28 &  !din_almost_full_7_29 &  !din_almost_full_7_30 &  !din_almost_full_7_31 &   1;
    //in_ready <= !in_eop; //create a gap
    
    in_data_r1 <= in_convt;
    in_data_r2 <= in_data_r1;

    //only valid when the input is dequeued. 
    in_valid_r1 <= in_valid;
    in_valid_r2 <= in_valid_r1;
    in_sop_r1 <= in_sop;
    in_sop_r2 <= in_sop_r1;
    in_eop_r1 <= in_eop;
    in_eop_r2 <= in_eop_r1;
    in_empty_r1 <= in_empty;
    in_empty_r2 <= in_empty_r1;
end

assign gap = (in_eop & in_valid & in_ready);

always@(posedge clk)begin
    if(rst)begin
        out_meta_valid <= 0;
    end else begin
        if(out_new_pkt)begin
            out_meta_valid <= 1;
        end else begin
            out_meta_valid <= 0;
        end
    end
    if(out_new_pkt)begin
        out_meta_data <= internal_meta_data;
        out_meta_data.pkt_flags <= PKT_DONE;
    end
end

assign internal_meta_ready = out_new_pkt;
//assign in_meta_ready = in_ready;

always@(posedge clk)begin
    din_valid_0_0 <= out_new_pkt | hash_out_valid_filter_0_0;
    din_valid_0_0_r1 <= din_valid_0_0;
    din_valid_0_0_r2 <= din_valid_0_0_r1;

    din_0_0.data <= hash_out_valid_filter_0_0 ? hash_out_0_0 : 0;
    din_0_0.last <= out_new_pkt;
    din_0_0.bucket <= 0;


    din_0_0_r1 <= din_0_0;
    din_0_0_r2 <= din_0_0_r1;
    din_valid_0_1 <= out_new_pkt | hash_out_valid_filter_0_1;
    din_valid_0_1_r1 <= din_valid_0_1;
    din_valid_0_1_r2 <= din_valid_0_1_r1;

    din_0_1.data <= hash_out_valid_filter_0_1 ? hash_out_0_1 : 0;
    din_0_1.last <= out_new_pkt;
    din_0_1.bucket <= 0;


    din_0_1_r1 <= din_0_1;
    din_0_1_r2 <= din_0_1_r1;
    din_valid_0_2 <= out_new_pkt | hash_out_valid_filter_0_2;
    din_valid_0_2_r1 <= din_valid_0_2;
    din_valid_0_2_r2 <= din_valid_0_2_r1;

    din_0_2.data <= hash_out_valid_filter_0_2 ? hash_out_0_2 : 0;
    din_0_2.last <= out_new_pkt;
    din_0_2.bucket <= 0;


    din_0_2_r1 <= din_0_2;
    din_0_2_r2 <= din_0_2_r1;
    din_valid_0_3 <= out_new_pkt | hash_out_valid_filter_0_3;
    din_valid_0_3_r1 <= din_valid_0_3;
    din_valid_0_3_r2 <= din_valid_0_3_r1;

    din_0_3.data <= hash_out_valid_filter_0_3 ? hash_out_0_3 : 0;
    din_0_3.last <= out_new_pkt;
    din_0_3.bucket <= 0;


    din_0_3_r1 <= din_0_3;
    din_0_3_r2 <= din_0_3_r1;
    din_valid_0_4 <= out_new_pkt | hash_out_valid_filter_0_4;
    din_valid_0_4_r1 <= din_valid_0_4;
    din_valid_0_4_r2 <= din_valid_0_4_r1;

    din_0_4.data <= hash_out_valid_filter_0_4 ? hash_out_0_4 : 0;
    din_0_4.last <= out_new_pkt;
    din_0_4.bucket <= 0;


    din_0_4_r1 <= din_0_4;
    din_0_4_r2 <= din_0_4_r1;
    din_valid_0_5 <= out_new_pkt | hash_out_valid_filter_0_5;
    din_valid_0_5_r1 <= din_valid_0_5;
    din_valid_0_5_r2 <= din_valid_0_5_r1;

    din_0_5.data <= hash_out_valid_filter_0_5 ? hash_out_0_5 : 0;
    din_0_5.last <= out_new_pkt;
    din_0_5.bucket <= 0;


    din_0_5_r1 <= din_0_5;
    din_0_5_r2 <= din_0_5_r1;
    din_valid_0_6 <= out_new_pkt | hash_out_valid_filter_0_6;
    din_valid_0_6_r1 <= din_valid_0_6;
    din_valid_0_6_r2 <= din_valid_0_6_r1;

    din_0_6.data <= hash_out_valid_filter_0_6 ? hash_out_0_6 : 0;
    din_0_6.last <= out_new_pkt;
    din_0_6.bucket <= 0;


    din_0_6_r1 <= din_0_6;
    din_0_6_r2 <= din_0_6_r1;
    din_valid_0_7 <= out_new_pkt | hash_out_valid_filter_0_7;
    din_valid_0_7_r1 <= din_valid_0_7;
    din_valid_0_7_r2 <= din_valid_0_7_r1;

    din_0_7.data <= hash_out_valid_filter_0_7 ? hash_out_0_7 : 0;
    din_0_7.last <= out_new_pkt;
    din_0_7.bucket <= 0;


    din_0_7_r1 <= din_0_7;
    din_0_7_r2 <= din_0_7_r1;
    din_valid_0_8 <= out_new_pkt | hash_out_valid_filter_0_8;
    din_valid_0_8_r1 <= din_valid_0_8;
    din_valid_0_8_r2 <= din_valid_0_8_r1;

    din_0_8.data <= hash_out_valid_filter_0_8 ? hash_out_0_8 : 0;
    din_0_8.last <= out_new_pkt;
    din_0_8.bucket <= 0;


    din_0_8_r1 <= din_0_8;
    din_0_8_r2 <= din_0_8_r1;
    din_valid_0_9 <= out_new_pkt | hash_out_valid_filter_0_9;
    din_valid_0_9_r1 <= din_valid_0_9;
    din_valid_0_9_r2 <= din_valid_0_9_r1;

    din_0_9.data <= hash_out_valid_filter_0_9 ? hash_out_0_9 : 0;
    din_0_9.last <= out_new_pkt;
    din_0_9.bucket <= 0;


    din_0_9_r1 <= din_0_9;
    din_0_9_r2 <= din_0_9_r1;
    din_valid_0_10 <= out_new_pkt | hash_out_valid_filter_0_10;
    din_valid_0_10_r1 <= din_valid_0_10;
    din_valid_0_10_r2 <= din_valid_0_10_r1;

    din_0_10.data <= hash_out_valid_filter_0_10 ? hash_out_0_10 : 0;
    din_0_10.last <= out_new_pkt;
    din_0_10.bucket <= 0;


    din_0_10_r1 <= din_0_10;
    din_0_10_r2 <= din_0_10_r1;
    din_valid_0_11 <= out_new_pkt | hash_out_valid_filter_0_11;
    din_valid_0_11_r1 <= din_valid_0_11;
    din_valid_0_11_r2 <= din_valid_0_11_r1;

    din_0_11.data <= hash_out_valid_filter_0_11 ? hash_out_0_11 : 0;
    din_0_11.last <= out_new_pkt;
    din_0_11.bucket <= 0;


    din_0_11_r1 <= din_0_11;
    din_0_11_r2 <= din_0_11_r1;
    din_valid_0_12 <= out_new_pkt | hash_out_valid_filter_0_12;
    din_valid_0_12_r1 <= din_valid_0_12;
    din_valid_0_12_r2 <= din_valid_0_12_r1;

    din_0_12.data <= hash_out_valid_filter_0_12 ? hash_out_0_12 : 0;
    din_0_12.last <= out_new_pkt;
    din_0_12.bucket <= 0;


    din_0_12_r1 <= din_0_12;
    din_0_12_r2 <= din_0_12_r1;
    din_valid_0_13 <= out_new_pkt | hash_out_valid_filter_0_13;
    din_valid_0_13_r1 <= din_valid_0_13;
    din_valid_0_13_r2 <= din_valid_0_13_r1;

    din_0_13.data <= hash_out_valid_filter_0_13 ? hash_out_0_13 : 0;
    din_0_13.last <= out_new_pkt;
    din_0_13.bucket <= 0;


    din_0_13_r1 <= din_0_13;
    din_0_13_r2 <= din_0_13_r1;
    din_valid_0_14 <= out_new_pkt | hash_out_valid_filter_0_14;
    din_valid_0_14_r1 <= din_valid_0_14;
    din_valid_0_14_r2 <= din_valid_0_14_r1;

    din_0_14.data <= hash_out_valid_filter_0_14 ? hash_out_0_14 : 0;
    din_0_14.last <= out_new_pkt;
    din_0_14.bucket <= 0;


    din_0_14_r1 <= din_0_14;
    din_0_14_r2 <= din_0_14_r1;
    din_valid_0_15 <= out_new_pkt | hash_out_valid_filter_0_15;
    din_valid_0_15_r1 <= din_valid_0_15;
    din_valid_0_15_r2 <= din_valid_0_15_r1;

    din_0_15.data <= hash_out_valid_filter_0_15 ? hash_out_0_15 : 0;
    din_0_15.last <= out_new_pkt;
    din_0_15.bucket <= 0;


    din_0_15_r1 <= din_0_15;
    din_0_15_r2 <= din_0_15_r1;
    din_valid_0_16 <= out_new_pkt | hash_out_valid_filter_0_16;
    din_valid_0_16_r1 <= din_valid_0_16;
    din_valid_0_16_r2 <= din_valid_0_16_r1;

    din_0_16.data <= hash_out_valid_filter_0_16 ? hash_out_0_16 : 0;
    din_0_16.last <= out_new_pkt;
    din_0_16.bucket <= 0;


    din_0_16_r1 <= din_0_16;
    din_0_16_r2 <= din_0_16_r1;
    din_valid_0_17 <= out_new_pkt | hash_out_valid_filter_0_17;
    din_valid_0_17_r1 <= din_valid_0_17;
    din_valid_0_17_r2 <= din_valid_0_17_r1;

    din_0_17.data <= hash_out_valid_filter_0_17 ? hash_out_0_17 : 0;
    din_0_17.last <= out_new_pkt;
    din_0_17.bucket <= 0;


    din_0_17_r1 <= din_0_17;
    din_0_17_r2 <= din_0_17_r1;
    din_valid_0_18 <= out_new_pkt | hash_out_valid_filter_0_18;
    din_valid_0_18_r1 <= din_valid_0_18;
    din_valid_0_18_r2 <= din_valid_0_18_r1;

    din_0_18.data <= hash_out_valid_filter_0_18 ? hash_out_0_18 : 0;
    din_0_18.last <= out_new_pkt;
    din_0_18.bucket <= 0;


    din_0_18_r1 <= din_0_18;
    din_0_18_r2 <= din_0_18_r1;
    din_valid_0_19 <= out_new_pkt | hash_out_valid_filter_0_19;
    din_valid_0_19_r1 <= din_valid_0_19;
    din_valid_0_19_r2 <= din_valid_0_19_r1;

    din_0_19.data <= hash_out_valid_filter_0_19 ? hash_out_0_19 : 0;
    din_0_19.last <= out_new_pkt;
    din_0_19.bucket <= 0;


    din_0_19_r1 <= din_0_19;
    din_0_19_r2 <= din_0_19_r1;
    din_valid_0_20 <= out_new_pkt | hash_out_valid_filter_0_20;
    din_valid_0_20_r1 <= din_valid_0_20;
    din_valid_0_20_r2 <= din_valid_0_20_r1;

    din_0_20.data <= hash_out_valid_filter_0_20 ? hash_out_0_20 : 0;
    din_0_20.last <= out_new_pkt;
    din_0_20.bucket <= 0;


    din_0_20_r1 <= din_0_20;
    din_0_20_r2 <= din_0_20_r1;
    din_valid_0_21 <= out_new_pkt | hash_out_valid_filter_0_21;
    din_valid_0_21_r1 <= din_valid_0_21;
    din_valid_0_21_r2 <= din_valid_0_21_r1;

    din_0_21.data <= hash_out_valid_filter_0_21 ? hash_out_0_21 : 0;
    din_0_21.last <= out_new_pkt;
    din_0_21.bucket <= 0;


    din_0_21_r1 <= din_0_21;
    din_0_21_r2 <= din_0_21_r1;
    din_valid_0_22 <= out_new_pkt | hash_out_valid_filter_0_22;
    din_valid_0_22_r1 <= din_valid_0_22;
    din_valid_0_22_r2 <= din_valid_0_22_r1;

    din_0_22.data <= hash_out_valid_filter_0_22 ? hash_out_0_22 : 0;
    din_0_22.last <= out_new_pkt;
    din_0_22.bucket <= 0;


    din_0_22_r1 <= din_0_22;
    din_0_22_r2 <= din_0_22_r1;
    din_valid_0_23 <= out_new_pkt | hash_out_valid_filter_0_23;
    din_valid_0_23_r1 <= din_valid_0_23;
    din_valid_0_23_r2 <= din_valid_0_23_r1;

    din_0_23.data <= hash_out_valid_filter_0_23 ? hash_out_0_23 : 0;
    din_0_23.last <= out_new_pkt;
    din_0_23.bucket <= 0;


    din_0_23_r1 <= din_0_23;
    din_0_23_r2 <= din_0_23_r1;
    din_valid_0_24 <= out_new_pkt | hash_out_valid_filter_0_24;
    din_valid_0_24_r1 <= din_valid_0_24;
    din_valid_0_24_r2 <= din_valid_0_24_r1;

    din_0_24.data <= hash_out_valid_filter_0_24 ? hash_out_0_24 : 0;
    din_0_24.last <= out_new_pkt;
    din_0_24.bucket <= 0;


    din_0_24_r1 <= din_0_24;
    din_0_24_r2 <= din_0_24_r1;
    din_valid_0_25 <= out_new_pkt | hash_out_valid_filter_0_25;
    din_valid_0_25_r1 <= din_valid_0_25;
    din_valid_0_25_r2 <= din_valid_0_25_r1;

    din_0_25.data <= hash_out_valid_filter_0_25 ? hash_out_0_25 : 0;
    din_0_25.last <= out_new_pkt;
    din_0_25.bucket <= 0;


    din_0_25_r1 <= din_0_25;
    din_0_25_r2 <= din_0_25_r1;
    din_valid_0_26 <= out_new_pkt | hash_out_valid_filter_0_26;
    din_valid_0_26_r1 <= din_valid_0_26;
    din_valid_0_26_r2 <= din_valid_0_26_r1;

    din_0_26.data <= hash_out_valid_filter_0_26 ? hash_out_0_26 : 0;
    din_0_26.last <= out_new_pkt;
    din_0_26.bucket <= 0;


    din_0_26_r1 <= din_0_26;
    din_0_26_r2 <= din_0_26_r1;
    din_valid_0_27 <= out_new_pkt | hash_out_valid_filter_0_27;
    din_valid_0_27_r1 <= din_valid_0_27;
    din_valid_0_27_r2 <= din_valid_0_27_r1;

    din_0_27.data <= hash_out_valid_filter_0_27 ? hash_out_0_27 : 0;
    din_0_27.last <= out_new_pkt;
    din_0_27.bucket <= 0;


    din_0_27_r1 <= din_0_27;
    din_0_27_r2 <= din_0_27_r1;
    din_valid_0_28 <= out_new_pkt | hash_out_valid_filter_0_28;
    din_valid_0_28_r1 <= din_valid_0_28;
    din_valid_0_28_r2 <= din_valid_0_28_r1;

    din_0_28.data <= hash_out_valid_filter_0_28 ? hash_out_0_28 : 0;
    din_0_28.last <= out_new_pkt;
    din_0_28.bucket <= 0;


    din_0_28_r1 <= din_0_28;
    din_0_28_r2 <= din_0_28_r1;
    din_valid_0_29 <= out_new_pkt | hash_out_valid_filter_0_29;
    din_valid_0_29_r1 <= din_valid_0_29;
    din_valid_0_29_r2 <= din_valid_0_29_r1;

    din_0_29.data <= hash_out_valid_filter_0_29 ? hash_out_0_29 : 0;
    din_0_29.last <= out_new_pkt;
    din_0_29.bucket <= 0;


    din_0_29_r1 <= din_0_29;
    din_0_29_r2 <= din_0_29_r1;
    din_valid_0_30 <= out_new_pkt | hash_out_valid_filter_0_30;
    din_valid_0_30_r1 <= din_valid_0_30;
    din_valid_0_30_r2 <= din_valid_0_30_r1;

    din_0_30.data <= hash_out_valid_filter_0_30 ? hash_out_0_30 : 0;
    din_0_30.last <= out_new_pkt;
    din_0_30.bucket <= 0;


    din_0_30_r1 <= din_0_30;
    din_0_30_r2 <= din_0_30_r1;
    din_valid_0_31 <= out_new_pkt | hash_out_valid_filter_0_31;
    din_valid_0_31_r1 <= din_valid_0_31;
    din_valid_0_31_r2 <= din_valid_0_31_r1;

    din_0_31.data <= hash_out_valid_filter_0_31 ? hash_out_0_31 : 0;
    din_0_31.last <= out_new_pkt;
    din_0_31.bucket <= 0;


    din_0_31_r1 <= din_0_31;
    din_0_31_r2 <= din_0_31_r1;
    din_valid_1_0 <= out_new_pkt | hash_out_valid_filter_1_0;
    din_valid_1_0_r1 <= din_valid_1_0;
    din_valid_1_0_r2 <= din_valid_1_0_r1;

    din_1_0.data <= hash_out_valid_filter_1_0 ? hash_out_1_0 : 0;
    din_1_0.last <= out_new_pkt;
    din_1_0.bucket <= 1;


    din_1_0_r1 <= din_1_0;
    din_1_0_r2 <= din_1_0_r1;
    din_valid_1_1 <= out_new_pkt | hash_out_valid_filter_1_1;
    din_valid_1_1_r1 <= din_valid_1_1;
    din_valid_1_1_r2 <= din_valid_1_1_r1;

    din_1_1.data <= hash_out_valid_filter_1_1 ? hash_out_1_1 : 0;
    din_1_1.last <= out_new_pkt;
    din_1_1.bucket <= 1;


    din_1_1_r1 <= din_1_1;
    din_1_1_r2 <= din_1_1_r1;
    din_valid_1_2 <= out_new_pkt | hash_out_valid_filter_1_2;
    din_valid_1_2_r1 <= din_valid_1_2;
    din_valid_1_2_r2 <= din_valid_1_2_r1;

    din_1_2.data <= hash_out_valid_filter_1_2 ? hash_out_1_2 : 0;
    din_1_2.last <= out_new_pkt;
    din_1_2.bucket <= 1;


    din_1_2_r1 <= din_1_2;
    din_1_2_r2 <= din_1_2_r1;
    din_valid_1_3 <= out_new_pkt | hash_out_valid_filter_1_3;
    din_valid_1_3_r1 <= din_valid_1_3;
    din_valid_1_3_r2 <= din_valid_1_3_r1;

    din_1_3.data <= hash_out_valid_filter_1_3 ? hash_out_1_3 : 0;
    din_1_3.last <= out_new_pkt;
    din_1_3.bucket <= 1;


    din_1_3_r1 <= din_1_3;
    din_1_3_r2 <= din_1_3_r1;
    din_valid_1_4 <= out_new_pkt | hash_out_valid_filter_1_4;
    din_valid_1_4_r1 <= din_valid_1_4;
    din_valid_1_4_r2 <= din_valid_1_4_r1;

    din_1_4.data <= hash_out_valid_filter_1_4 ? hash_out_1_4 : 0;
    din_1_4.last <= out_new_pkt;
    din_1_4.bucket <= 1;


    din_1_4_r1 <= din_1_4;
    din_1_4_r2 <= din_1_4_r1;
    din_valid_1_5 <= out_new_pkt | hash_out_valid_filter_1_5;
    din_valid_1_5_r1 <= din_valid_1_5;
    din_valid_1_5_r2 <= din_valid_1_5_r1;

    din_1_5.data <= hash_out_valid_filter_1_5 ? hash_out_1_5 : 0;
    din_1_5.last <= out_new_pkt;
    din_1_5.bucket <= 1;


    din_1_5_r1 <= din_1_5;
    din_1_5_r2 <= din_1_5_r1;
    din_valid_1_6 <= out_new_pkt | hash_out_valid_filter_1_6;
    din_valid_1_6_r1 <= din_valid_1_6;
    din_valid_1_6_r2 <= din_valid_1_6_r1;

    din_1_6.data <= hash_out_valid_filter_1_6 ? hash_out_1_6 : 0;
    din_1_6.last <= out_new_pkt;
    din_1_6.bucket <= 1;


    din_1_6_r1 <= din_1_6;
    din_1_6_r2 <= din_1_6_r1;
    din_valid_1_7 <= out_new_pkt | hash_out_valid_filter_1_7;
    din_valid_1_7_r1 <= din_valid_1_7;
    din_valid_1_7_r2 <= din_valid_1_7_r1;

    din_1_7.data <= hash_out_valid_filter_1_7 ? hash_out_1_7 : 0;
    din_1_7.last <= out_new_pkt;
    din_1_7.bucket <= 1;


    din_1_7_r1 <= din_1_7;
    din_1_7_r2 <= din_1_7_r1;
    din_valid_1_8 <= out_new_pkt | hash_out_valid_filter_1_8;
    din_valid_1_8_r1 <= din_valid_1_8;
    din_valid_1_8_r2 <= din_valid_1_8_r1;

    din_1_8.data <= hash_out_valid_filter_1_8 ? hash_out_1_8 : 0;
    din_1_8.last <= out_new_pkt;
    din_1_8.bucket <= 1;


    din_1_8_r1 <= din_1_8;
    din_1_8_r2 <= din_1_8_r1;
    din_valid_1_9 <= out_new_pkt | hash_out_valid_filter_1_9;
    din_valid_1_9_r1 <= din_valid_1_9;
    din_valid_1_9_r2 <= din_valid_1_9_r1;

    din_1_9.data <= hash_out_valid_filter_1_9 ? hash_out_1_9 : 0;
    din_1_9.last <= out_new_pkt;
    din_1_9.bucket <= 1;


    din_1_9_r1 <= din_1_9;
    din_1_9_r2 <= din_1_9_r1;
    din_valid_1_10 <= out_new_pkt | hash_out_valid_filter_1_10;
    din_valid_1_10_r1 <= din_valid_1_10;
    din_valid_1_10_r2 <= din_valid_1_10_r1;

    din_1_10.data <= hash_out_valid_filter_1_10 ? hash_out_1_10 : 0;
    din_1_10.last <= out_new_pkt;
    din_1_10.bucket <= 1;


    din_1_10_r1 <= din_1_10;
    din_1_10_r2 <= din_1_10_r1;
    din_valid_1_11 <= out_new_pkt | hash_out_valid_filter_1_11;
    din_valid_1_11_r1 <= din_valid_1_11;
    din_valid_1_11_r2 <= din_valid_1_11_r1;

    din_1_11.data <= hash_out_valid_filter_1_11 ? hash_out_1_11 : 0;
    din_1_11.last <= out_new_pkt;
    din_1_11.bucket <= 1;


    din_1_11_r1 <= din_1_11;
    din_1_11_r2 <= din_1_11_r1;
    din_valid_1_12 <= out_new_pkt | hash_out_valid_filter_1_12;
    din_valid_1_12_r1 <= din_valid_1_12;
    din_valid_1_12_r2 <= din_valid_1_12_r1;

    din_1_12.data <= hash_out_valid_filter_1_12 ? hash_out_1_12 : 0;
    din_1_12.last <= out_new_pkt;
    din_1_12.bucket <= 1;


    din_1_12_r1 <= din_1_12;
    din_1_12_r2 <= din_1_12_r1;
    din_valid_1_13 <= out_new_pkt | hash_out_valid_filter_1_13;
    din_valid_1_13_r1 <= din_valid_1_13;
    din_valid_1_13_r2 <= din_valid_1_13_r1;

    din_1_13.data <= hash_out_valid_filter_1_13 ? hash_out_1_13 : 0;
    din_1_13.last <= out_new_pkt;
    din_1_13.bucket <= 1;


    din_1_13_r1 <= din_1_13;
    din_1_13_r2 <= din_1_13_r1;
    din_valid_1_14 <= out_new_pkt | hash_out_valid_filter_1_14;
    din_valid_1_14_r1 <= din_valid_1_14;
    din_valid_1_14_r2 <= din_valid_1_14_r1;

    din_1_14.data <= hash_out_valid_filter_1_14 ? hash_out_1_14 : 0;
    din_1_14.last <= out_new_pkt;
    din_1_14.bucket <= 1;


    din_1_14_r1 <= din_1_14;
    din_1_14_r2 <= din_1_14_r1;
    din_valid_1_15 <= out_new_pkt | hash_out_valid_filter_1_15;
    din_valid_1_15_r1 <= din_valid_1_15;
    din_valid_1_15_r2 <= din_valid_1_15_r1;

    din_1_15.data <= hash_out_valid_filter_1_15 ? hash_out_1_15 : 0;
    din_1_15.last <= out_new_pkt;
    din_1_15.bucket <= 1;


    din_1_15_r1 <= din_1_15;
    din_1_15_r2 <= din_1_15_r1;
    din_valid_1_16 <= out_new_pkt | hash_out_valid_filter_1_16;
    din_valid_1_16_r1 <= din_valid_1_16;
    din_valid_1_16_r2 <= din_valid_1_16_r1;

    din_1_16.data <= hash_out_valid_filter_1_16 ? hash_out_1_16 : 0;
    din_1_16.last <= out_new_pkt;
    din_1_16.bucket <= 1;


    din_1_16_r1 <= din_1_16;
    din_1_16_r2 <= din_1_16_r1;
    din_valid_1_17 <= out_new_pkt | hash_out_valid_filter_1_17;
    din_valid_1_17_r1 <= din_valid_1_17;
    din_valid_1_17_r2 <= din_valid_1_17_r1;

    din_1_17.data <= hash_out_valid_filter_1_17 ? hash_out_1_17 : 0;
    din_1_17.last <= out_new_pkt;
    din_1_17.bucket <= 1;


    din_1_17_r1 <= din_1_17;
    din_1_17_r2 <= din_1_17_r1;
    din_valid_1_18 <= out_new_pkt | hash_out_valid_filter_1_18;
    din_valid_1_18_r1 <= din_valid_1_18;
    din_valid_1_18_r2 <= din_valid_1_18_r1;

    din_1_18.data <= hash_out_valid_filter_1_18 ? hash_out_1_18 : 0;
    din_1_18.last <= out_new_pkt;
    din_1_18.bucket <= 1;


    din_1_18_r1 <= din_1_18;
    din_1_18_r2 <= din_1_18_r1;
    din_valid_1_19 <= out_new_pkt | hash_out_valid_filter_1_19;
    din_valid_1_19_r1 <= din_valid_1_19;
    din_valid_1_19_r2 <= din_valid_1_19_r1;

    din_1_19.data <= hash_out_valid_filter_1_19 ? hash_out_1_19 : 0;
    din_1_19.last <= out_new_pkt;
    din_1_19.bucket <= 1;


    din_1_19_r1 <= din_1_19;
    din_1_19_r2 <= din_1_19_r1;
    din_valid_1_20 <= out_new_pkt | hash_out_valid_filter_1_20;
    din_valid_1_20_r1 <= din_valid_1_20;
    din_valid_1_20_r2 <= din_valid_1_20_r1;

    din_1_20.data <= hash_out_valid_filter_1_20 ? hash_out_1_20 : 0;
    din_1_20.last <= out_new_pkt;
    din_1_20.bucket <= 1;


    din_1_20_r1 <= din_1_20;
    din_1_20_r2 <= din_1_20_r1;
    din_valid_1_21 <= out_new_pkt | hash_out_valid_filter_1_21;
    din_valid_1_21_r1 <= din_valid_1_21;
    din_valid_1_21_r2 <= din_valid_1_21_r1;

    din_1_21.data <= hash_out_valid_filter_1_21 ? hash_out_1_21 : 0;
    din_1_21.last <= out_new_pkt;
    din_1_21.bucket <= 1;


    din_1_21_r1 <= din_1_21;
    din_1_21_r2 <= din_1_21_r1;
    din_valid_1_22 <= out_new_pkt | hash_out_valid_filter_1_22;
    din_valid_1_22_r1 <= din_valid_1_22;
    din_valid_1_22_r2 <= din_valid_1_22_r1;

    din_1_22.data <= hash_out_valid_filter_1_22 ? hash_out_1_22 : 0;
    din_1_22.last <= out_new_pkt;
    din_1_22.bucket <= 1;


    din_1_22_r1 <= din_1_22;
    din_1_22_r2 <= din_1_22_r1;
    din_valid_1_23 <= out_new_pkt | hash_out_valid_filter_1_23;
    din_valid_1_23_r1 <= din_valid_1_23;
    din_valid_1_23_r2 <= din_valid_1_23_r1;

    din_1_23.data <= hash_out_valid_filter_1_23 ? hash_out_1_23 : 0;
    din_1_23.last <= out_new_pkt;
    din_1_23.bucket <= 1;


    din_1_23_r1 <= din_1_23;
    din_1_23_r2 <= din_1_23_r1;
    din_valid_1_24 <= out_new_pkt | hash_out_valid_filter_1_24;
    din_valid_1_24_r1 <= din_valid_1_24;
    din_valid_1_24_r2 <= din_valid_1_24_r1;

    din_1_24.data <= hash_out_valid_filter_1_24 ? hash_out_1_24 : 0;
    din_1_24.last <= out_new_pkt;
    din_1_24.bucket <= 1;


    din_1_24_r1 <= din_1_24;
    din_1_24_r2 <= din_1_24_r1;
    din_valid_1_25 <= out_new_pkt | hash_out_valid_filter_1_25;
    din_valid_1_25_r1 <= din_valid_1_25;
    din_valid_1_25_r2 <= din_valid_1_25_r1;

    din_1_25.data <= hash_out_valid_filter_1_25 ? hash_out_1_25 : 0;
    din_1_25.last <= out_new_pkt;
    din_1_25.bucket <= 1;


    din_1_25_r1 <= din_1_25;
    din_1_25_r2 <= din_1_25_r1;
    din_valid_1_26 <= out_new_pkt | hash_out_valid_filter_1_26;
    din_valid_1_26_r1 <= din_valid_1_26;
    din_valid_1_26_r2 <= din_valid_1_26_r1;

    din_1_26.data <= hash_out_valid_filter_1_26 ? hash_out_1_26 : 0;
    din_1_26.last <= out_new_pkt;
    din_1_26.bucket <= 1;


    din_1_26_r1 <= din_1_26;
    din_1_26_r2 <= din_1_26_r1;
    din_valid_1_27 <= out_new_pkt | hash_out_valid_filter_1_27;
    din_valid_1_27_r1 <= din_valid_1_27;
    din_valid_1_27_r2 <= din_valid_1_27_r1;

    din_1_27.data <= hash_out_valid_filter_1_27 ? hash_out_1_27 : 0;
    din_1_27.last <= out_new_pkt;
    din_1_27.bucket <= 1;


    din_1_27_r1 <= din_1_27;
    din_1_27_r2 <= din_1_27_r1;
    din_valid_1_28 <= out_new_pkt | hash_out_valid_filter_1_28;
    din_valid_1_28_r1 <= din_valid_1_28;
    din_valid_1_28_r2 <= din_valid_1_28_r1;

    din_1_28.data <= hash_out_valid_filter_1_28 ? hash_out_1_28 : 0;
    din_1_28.last <= out_new_pkt;
    din_1_28.bucket <= 1;


    din_1_28_r1 <= din_1_28;
    din_1_28_r2 <= din_1_28_r1;
    din_valid_1_29 <= out_new_pkt | hash_out_valid_filter_1_29;
    din_valid_1_29_r1 <= din_valid_1_29;
    din_valid_1_29_r2 <= din_valid_1_29_r1;

    din_1_29.data <= hash_out_valid_filter_1_29 ? hash_out_1_29 : 0;
    din_1_29.last <= out_new_pkt;
    din_1_29.bucket <= 1;


    din_1_29_r1 <= din_1_29;
    din_1_29_r2 <= din_1_29_r1;
    din_valid_1_30 <= out_new_pkt | hash_out_valid_filter_1_30;
    din_valid_1_30_r1 <= din_valid_1_30;
    din_valid_1_30_r2 <= din_valid_1_30_r1;

    din_1_30.data <= hash_out_valid_filter_1_30 ? hash_out_1_30 : 0;
    din_1_30.last <= out_new_pkt;
    din_1_30.bucket <= 1;


    din_1_30_r1 <= din_1_30;
    din_1_30_r2 <= din_1_30_r1;
    din_valid_1_31 <= out_new_pkt | hash_out_valid_filter_1_31;
    din_valid_1_31_r1 <= din_valid_1_31;
    din_valid_1_31_r2 <= din_valid_1_31_r1;

    din_1_31.data <= hash_out_valid_filter_1_31 ? hash_out_1_31 : 0;
    din_1_31.last <= out_new_pkt;
    din_1_31.bucket <= 1;


    din_1_31_r1 <= din_1_31;
    din_1_31_r2 <= din_1_31_r1;
    din_valid_2_0 <= out_new_pkt | hash_out_valid_filter_2_0;
    din_valid_2_0_r1 <= din_valid_2_0;
    din_valid_2_0_r2 <= din_valid_2_0_r1;

    din_2_0.data <= hash_out_valid_filter_2_0 ? hash_out_2_0 : 0;
    din_2_0.last <= out_new_pkt;
    din_2_0.bucket <= 2;


    din_2_0_r1 <= din_2_0;
    din_2_0_r2 <= din_2_0_r1;
    din_valid_2_1 <= out_new_pkt | hash_out_valid_filter_2_1;
    din_valid_2_1_r1 <= din_valid_2_1;
    din_valid_2_1_r2 <= din_valid_2_1_r1;

    din_2_1.data <= hash_out_valid_filter_2_1 ? hash_out_2_1 : 0;
    din_2_1.last <= out_new_pkt;
    din_2_1.bucket <= 2;


    din_2_1_r1 <= din_2_1;
    din_2_1_r2 <= din_2_1_r1;
    din_valid_2_2 <= out_new_pkt | hash_out_valid_filter_2_2;
    din_valid_2_2_r1 <= din_valid_2_2;
    din_valid_2_2_r2 <= din_valid_2_2_r1;

    din_2_2.data <= hash_out_valid_filter_2_2 ? hash_out_2_2 : 0;
    din_2_2.last <= out_new_pkt;
    din_2_2.bucket <= 2;


    din_2_2_r1 <= din_2_2;
    din_2_2_r2 <= din_2_2_r1;
    din_valid_2_3 <= out_new_pkt | hash_out_valid_filter_2_3;
    din_valid_2_3_r1 <= din_valid_2_3;
    din_valid_2_3_r2 <= din_valid_2_3_r1;

    din_2_3.data <= hash_out_valid_filter_2_3 ? hash_out_2_3 : 0;
    din_2_3.last <= out_new_pkt;
    din_2_3.bucket <= 2;


    din_2_3_r1 <= din_2_3;
    din_2_3_r2 <= din_2_3_r1;
    din_valid_2_4 <= out_new_pkt | hash_out_valid_filter_2_4;
    din_valid_2_4_r1 <= din_valid_2_4;
    din_valid_2_4_r2 <= din_valid_2_4_r1;

    din_2_4.data <= hash_out_valid_filter_2_4 ? hash_out_2_4 : 0;
    din_2_4.last <= out_new_pkt;
    din_2_4.bucket <= 2;


    din_2_4_r1 <= din_2_4;
    din_2_4_r2 <= din_2_4_r1;
    din_valid_2_5 <= out_new_pkt | hash_out_valid_filter_2_5;
    din_valid_2_5_r1 <= din_valid_2_5;
    din_valid_2_5_r2 <= din_valid_2_5_r1;

    din_2_5.data <= hash_out_valid_filter_2_5 ? hash_out_2_5 : 0;
    din_2_5.last <= out_new_pkt;
    din_2_5.bucket <= 2;


    din_2_5_r1 <= din_2_5;
    din_2_5_r2 <= din_2_5_r1;
    din_valid_2_6 <= out_new_pkt | hash_out_valid_filter_2_6;
    din_valid_2_6_r1 <= din_valid_2_6;
    din_valid_2_6_r2 <= din_valid_2_6_r1;

    din_2_6.data <= hash_out_valid_filter_2_6 ? hash_out_2_6 : 0;
    din_2_6.last <= out_new_pkt;
    din_2_6.bucket <= 2;


    din_2_6_r1 <= din_2_6;
    din_2_6_r2 <= din_2_6_r1;
    din_valid_2_7 <= out_new_pkt | hash_out_valid_filter_2_7;
    din_valid_2_7_r1 <= din_valid_2_7;
    din_valid_2_7_r2 <= din_valid_2_7_r1;

    din_2_7.data <= hash_out_valid_filter_2_7 ? hash_out_2_7 : 0;
    din_2_7.last <= out_new_pkt;
    din_2_7.bucket <= 2;


    din_2_7_r1 <= din_2_7;
    din_2_7_r2 <= din_2_7_r1;
    din_valid_2_8 <= out_new_pkt | hash_out_valid_filter_2_8;
    din_valid_2_8_r1 <= din_valid_2_8;
    din_valid_2_8_r2 <= din_valid_2_8_r1;

    din_2_8.data <= hash_out_valid_filter_2_8 ? hash_out_2_8 : 0;
    din_2_8.last <= out_new_pkt;
    din_2_8.bucket <= 2;


    din_2_8_r1 <= din_2_8;
    din_2_8_r2 <= din_2_8_r1;
    din_valid_2_9 <= out_new_pkt | hash_out_valid_filter_2_9;
    din_valid_2_9_r1 <= din_valid_2_9;
    din_valid_2_9_r2 <= din_valid_2_9_r1;

    din_2_9.data <= hash_out_valid_filter_2_9 ? hash_out_2_9 : 0;
    din_2_9.last <= out_new_pkt;
    din_2_9.bucket <= 2;


    din_2_9_r1 <= din_2_9;
    din_2_9_r2 <= din_2_9_r1;
    din_valid_2_10 <= out_new_pkt | hash_out_valid_filter_2_10;
    din_valid_2_10_r1 <= din_valid_2_10;
    din_valid_2_10_r2 <= din_valid_2_10_r1;

    din_2_10.data <= hash_out_valid_filter_2_10 ? hash_out_2_10 : 0;
    din_2_10.last <= out_new_pkt;
    din_2_10.bucket <= 2;


    din_2_10_r1 <= din_2_10;
    din_2_10_r2 <= din_2_10_r1;
    din_valid_2_11 <= out_new_pkt | hash_out_valid_filter_2_11;
    din_valid_2_11_r1 <= din_valid_2_11;
    din_valid_2_11_r2 <= din_valid_2_11_r1;

    din_2_11.data <= hash_out_valid_filter_2_11 ? hash_out_2_11 : 0;
    din_2_11.last <= out_new_pkt;
    din_2_11.bucket <= 2;


    din_2_11_r1 <= din_2_11;
    din_2_11_r2 <= din_2_11_r1;
    din_valid_2_12 <= out_new_pkt | hash_out_valid_filter_2_12;
    din_valid_2_12_r1 <= din_valid_2_12;
    din_valid_2_12_r2 <= din_valid_2_12_r1;

    din_2_12.data <= hash_out_valid_filter_2_12 ? hash_out_2_12 : 0;
    din_2_12.last <= out_new_pkt;
    din_2_12.bucket <= 2;


    din_2_12_r1 <= din_2_12;
    din_2_12_r2 <= din_2_12_r1;
    din_valid_2_13 <= out_new_pkt | hash_out_valid_filter_2_13;
    din_valid_2_13_r1 <= din_valid_2_13;
    din_valid_2_13_r2 <= din_valid_2_13_r1;

    din_2_13.data <= hash_out_valid_filter_2_13 ? hash_out_2_13 : 0;
    din_2_13.last <= out_new_pkt;
    din_2_13.bucket <= 2;


    din_2_13_r1 <= din_2_13;
    din_2_13_r2 <= din_2_13_r1;
    din_valid_2_14 <= out_new_pkt | hash_out_valid_filter_2_14;
    din_valid_2_14_r1 <= din_valid_2_14;
    din_valid_2_14_r2 <= din_valid_2_14_r1;

    din_2_14.data <= hash_out_valid_filter_2_14 ? hash_out_2_14 : 0;
    din_2_14.last <= out_new_pkt;
    din_2_14.bucket <= 2;


    din_2_14_r1 <= din_2_14;
    din_2_14_r2 <= din_2_14_r1;
    din_valid_2_15 <= out_new_pkt | hash_out_valid_filter_2_15;
    din_valid_2_15_r1 <= din_valid_2_15;
    din_valid_2_15_r2 <= din_valid_2_15_r1;

    din_2_15.data <= hash_out_valid_filter_2_15 ? hash_out_2_15 : 0;
    din_2_15.last <= out_new_pkt;
    din_2_15.bucket <= 2;


    din_2_15_r1 <= din_2_15;
    din_2_15_r2 <= din_2_15_r1;
    din_valid_2_16 <= out_new_pkt | hash_out_valid_filter_2_16;
    din_valid_2_16_r1 <= din_valid_2_16;
    din_valid_2_16_r2 <= din_valid_2_16_r1;

    din_2_16.data <= hash_out_valid_filter_2_16 ? hash_out_2_16 : 0;
    din_2_16.last <= out_new_pkt;
    din_2_16.bucket <= 2;


    din_2_16_r1 <= din_2_16;
    din_2_16_r2 <= din_2_16_r1;
    din_valid_2_17 <= out_new_pkt | hash_out_valid_filter_2_17;
    din_valid_2_17_r1 <= din_valid_2_17;
    din_valid_2_17_r2 <= din_valid_2_17_r1;

    din_2_17.data <= hash_out_valid_filter_2_17 ? hash_out_2_17 : 0;
    din_2_17.last <= out_new_pkt;
    din_2_17.bucket <= 2;


    din_2_17_r1 <= din_2_17;
    din_2_17_r2 <= din_2_17_r1;
    din_valid_2_18 <= out_new_pkt | hash_out_valid_filter_2_18;
    din_valid_2_18_r1 <= din_valid_2_18;
    din_valid_2_18_r2 <= din_valid_2_18_r1;

    din_2_18.data <= hash_out_valid_filter_2_18 ? hash_out_2_18 : 0;
    din_2_18.last <= out_new_pkt;
    din_2_18.bucket <= 2;


    din_2_18_r1 <= din_2_18;
    din_2_18_r2 <= din_2_18_r1;
    din_valid_2_19 <= out_new_pkt | hash_out_valid_filter_2_19;
    din_valid_2_19_r1 <= din_valid_2_19;
    din_valid_2_19_r2 <= din_valid_2_19_r1;

    din_2_19.data <= hash_out_valid_filter_2_19 ? hash_out_2_19 : 0;
    din_2_19.last <= out_new_pkt;
    din_2_19.bucket <= 2;


    din_2_19_r1 <= din_2_19;
    din_2_19_r2 <= din_2_19_r1;
    din_valid_2_20 <= out_new_pkt | hash_out_valid_filter_2_20;
    din_valid_2_20_r1 <= din_valid_2_20;
    din_valid_2_20_r2 <= din_valid_2_20_r1;

    din_2_20.data <= hash_out_valid_filter_2_20 ? hash_out_2_20 : 0;
    din_2_20.last <= out_new_pkt;
    din_2_20.bucket <= 2;


    din_2_20_r1 <= din_2_20;
    din_2_20_r2 <= din_2_20_r1;
    din_valid_2_21 <= out_new_pkt | hash_out_valid_filter_2_21;
    din_valid_2_21_r1 <= din_valid_2_21;
    din_valid_2_21_r2 <= din_valid_2_21_r1;

    din_2_21.data <= hash_out_valid_filter_2_21 ? hash_out_2_21 : 0;
    din_2_21.last <= out_new_pkt;
    din_2_21.bucket <= 2;


    din_2_21_r1 <= din_2_21;
    din_2_21_r2 <= din_2_21_r1;
    din_valid_2_22 <= out_new_pkt | hash_out_valid_filter_2_22;
    din_valid_2_22_r1 <= din_valid_2_22;
    din_valid_2_22_r2 <= din_valid_2_22_r1;

    din_2_22.data <= hash_out_valid_filter_2_22 ? hash_out_2_22 : 0;
    din_2_22.last <= out_new_pkt;
    din_2_22.bucket <= 2;


    din_2_22_r1 <= din_2_22;
    din_2_22_r2 <= din_2_22_r1;
    din_valid_2_23 <= out_new_pkt | hash_out_valid_filter_2_23;
    din_valid_2_23_r1 <= din_valid_2_23;
    din_valid_2_23_r2 <= din_valid_2_23_r1;

    din_2_23.data <= hash_out_valid_filter_2_23 ? hash_out_2_23 : 0;
    din_2_23.last <= out_new_pkt;
    din_2_23.bucket <= 2;


    din_2_23_r1 <= din_2_23;
    din_2_23_r2 <= din_2_23_r1;
    din_valid_2_24 <= out_new_pkt | hash_out_valid_filter_2_24;
    din_valid_2_24_r1 <= din_valid_2_24;
    din_valid_2_24_r2 <= din_valid_2_24_r1;

    din_2_24.data <= hash_out_valid_filter_2_24 ? hash_out_2_24 : 0;
    din_2_24.last <= out_new_pkt;
    din_2_24.bucket <= 2;


    din_2_24_r1 <= din_2_24;
    din_2_24_r2 <= din_2_24_r1;
    din_valid_2_25 <= out_new_pkt | hash_out_valid_filter_2_25;
    din_valid_2_25_r1 <= din_valid_2_25;
    din_valid_2_25_r2 <= din_valid_2_25_r1;

    din_2_25.data <= hash_out_valid_filter_2_25 ? hash_out_2_25 : 0;
    din_2_25.last <= out_new_pkt;
    din_2_25.bucket <= 2;


    din_2_25_r1 <= din_2_25;
    din_2_25_r2 <= din_2_25_r1;
    din_valid_2_26 <= out_new_pkt | hash_out_valid_filter_2_26;
    din_valid_2_26_r1 <= din_valid_2_26;
    din_valid_2_26_r2 <= din_valid_2_26_r1;

    din_2_26.data <= hash_out_valid_filter_2_26 ? hash_out_2_26 : 0;
    din_2_26.last <= out_new_pkt;
    din_2_26.bucket <= 2;


    din_2_26_r1 <= din_2_26;
    din_2_26_r2 <= din_2_26_r1;
    din_valid_2_27 <= out_new_pkt | hash_out_valid_filter_2_27;
    din_valid_2_27_r1 <= din_valid_2_27;
    din_valid_2_27_r2 <= din_valid_2_27_r1;

    din_2_27.data <= hash_out_valid_filter_2_27 ? hash_out_2_27 : 0;
    din_2_27.last <= out_new_pkt;
    din_2_27.bucket <= 2;


    din_2_27_r1 <= din_2_27;
    din_2_27_r2 <= din_2_27_r1;
    din_valid_2_28 <= out_new_pkt | hash_out_valid_filter_2_28;
    din_valid_2_28_r1 <= din_valid_2_28;
    din_valid_2_28_r2 <= din_valid_2_28_r1;

    din_2_28.data <= hash_out_valid_filter_2_28 ? hash_out_2_28 : 0;
    din_2_28.last <= out_new_pkt;
    din_2_28.bucket <= 2;


    din_2_28_r1 <= din_2_28;
    din_2_28_r2 <= din_2_28_r1;
    din_valid_2_29 <= out_new_pkt | hash_out_valid_filter_2_29;
    din_valid_2_29_r1 <= din_valid_2_29;
    din_valid_2_29_r2 <= din_valid_2_29_r1;

    din_2_29.data <= hash_out_valid_filter_2_29 ? hash_out_2_29 : 0;
    din_2_29.last <= out_new_pkt;
    din_2_29.bucket <= 2;


    din_2_29_r1 <= din_2_29;
    din_2_29_r2 <= din_2_29_r1;
    din_valid_2_30 <= out_new_pkt | hash_out_valid_filter_2_30;
    din_valid_2_30_r1 <= din_valid_2_30;
    din_valid_2_30_r2 <= din_valid_2_30_r1;

    din_2_30.data <= hash_out_valid_filter_2_30 ? hash_out_2_30 : 0;
    din_2_30.last <= out_new_pkt;
    din_2_30.bucket <= 2;


    din_2_30_r1 <= din_2_30;
    din_2_30_r2 <= din_2_30_r1;
    din_valid_2_31 <= out_new_pkt | hash_out_valid_filter_2_31;
    din_valid_2_31_r1 <= din_valid_2_31;
    din_valid_2_31_r2 <= din_valid_2_31_r1;

    din_2_31.data <= hash_out_valid_filter_2_31 ? hash_out_2_31 : 0;
    din_2_31.last <= out_new_pkt;
    din_2_31.bucket <= 2;


    din_2_31_r1 <= din_2_31;
    din_2_31_r2 <= din_2_31_r1;
    din_valid_3_0 <= out_new_pkt | hash_out_valid_filter_3_0;
    din_valid_3_0_r1 <= din_valid_3_0;
    din_valid_3_0_r2 <= din_valid_3_0_r1;

    din_3_0.data <= hash_out_valid_filter_3_0 ? hash_out_3_0 : 0;
    din_3_0.last <= out_new_pkt;
    din_3_0.bucket <= 3;


    din_3_0_r1 <= din_3_0;
    din_3_0_r2 <= din_3_0_r1;
    din_valid_3_1 <= out_new_pkt | hash_out_valid_filter_3_1;
    din_valid_3_1_r1 <= din_valid_3_1;
    din_valid_3_1_r2 <= din_valid_3_1_r1;

    din_3_1.data <= hash_out_valid_filter_3_1 ? hash_out_3_1 : 0;
    din_3_1.last <= out_new_pkt;
    din_3_1.bucket <= 3;


    din_3_1_r1 <= din_3_1;
    din_3_1_r2 <= din_3_1_r1;
    din_valid_3_2 <= out_new_pkt | hash_out_valid_filter_3_2;
    din_valid_3_2_r1 <= din_valid_3_2;
    din_valid_3_2_r2 <= din_valid_3_2_r1;

    din_3_2.data <= hash_out_valid_filter_3_2 ? hash_out_3_2 : 0;
    din_3_2.last <= out_new_pkt;
    din_3_2.bucket <= 3;


    din_3_2_r1 <= din_3_2;
    din_3_2_r2 <= din_3_2_r1;
    din_valid_3_3 <= out_new_pkt | hash_out_valid_filter_3_3;
    din_valid_3_3_r1 <= din_valid_3_3;
    din_valid_3_3_r2 <= din_valid_3_3_r1;

    din_3_3.data <= hash_out_valid_filter_3_3 ? hash_out_3_3 : 0;
    din_3_3.last <= out_new_pkt;
    din_3_3.bucket <= 3;


    din_3_3_r1 <= din_3_3;
    din_3_3_r2 <= din_3_3_r1;
    din_valid_3_4 <= out_new_pkt | hash_out_valid_filter_3_4;
    din_valid_3_4_r1 <= din_valid_3_4;
    din_valid_3_4_r2 <= din_valid_3_4_r1;

    din_3_4.data <= hash_out_valid_filter_3_4 ? hash_out_3_4 : 0;
    din_3_4.last <= out_new_pkt;
    din_3_4.bucket <= 3;


    din_3_4_r1 <= din_3_4;
    din_3_4_r2 <= din_3_4_r1;
    din_valid_3_5 <= out_new_pkt | hash_out_valid_filter_3_5;
    din_valid_3_5_r1 <= din_valid_3_5;
    din_valid_3_5_r2 <= din_valid_3_5_r1;

    din_3_5.data <= hash_out_valid_filter_3_5 ? hash_out_3_5 : 0;
    din_3_5.last <= out_new_pkt;
    din_3_5.bucket <= 3;


    din_3_5_r1 <= din_3_5;
    din_3_5_r2 <= din_3_5_r1;
    din_valid_3_6 <= out_new_pkt | hash_out_valid_filter_3_6;
    din_valid_3_6_r1 <= din_valid_3_6;
    din_valid_3_6_r2 <= din_valid_3_6_r1;

    din_3_6.data <= hash_out_valid_filter_3_6 ? hash_out_3_6 : 0;
    din_3_6.last <= out_new_pkt;
    din_3_6.bucket <= 3;


    din_3_6_r1 <= din_3_6;
    din_3_6_r2 <= din_3_6_r1;
    din_valid_3_7 <= out_new_pkt | hash_out_valid_filter_3_7;
    din_valid_3_7_r1 <= din_valid_3_7;
    din_valid_3_7_r2 <= din_valid_3_7_r1;

    din_3_7.data <= hash_out_valid_filter_3_7 ? hash_out_3_7 : 0;
    din_3_7.last <= out_new_pkt;
    din_3_7.bucket <= 3;


    din_3_7_r1 <= din_3_7;
    din_3_7_r2 <= din_3_7_r1;
    din_valid_3_8 <= out_new_pkt | hash_out_valid_filter_3_8;
    din_valid_3_8_r1 <= din_valid_3_8;
    din_valid_3_8_r2 <= din_valid_3_8_r1;

    din_3_8.data <= hash_out_valid_filter_3_8 ? hash_out_3_8 : 0;
    din_3_8.last <= out_new_pkt;
    din_3_8.bucket <= 3;


    din_3_8_r1 <= din_3_8;
    din_3_8_r2 <= din_3_8_r1;
    din_valid_3_9 <= out_new_pkt | hash_out_valid_filter_3_9;
    din_valid_3_9_r1 <= din_valid_3_9;
    din_valid_3_9_r2 <= din_valid_3_9_r1;

    din_3_9.data <= hash_out_valid_filter_3_9 ? hash_out_3_9 : 0;
    din_3_9.last <= out_new_pkt;
    din_3_9.bucket <= 3;


    din_3_9_r1 <= din_3_9;
    din_3_9_r2 <= din_3_9_r1;
    din_valid_3_10 <= out_new_pkt | hash_out_valid_filter_3_10;
    din_valid_3_10_r1 <= din_valid_3_10;
    din_valid_3_10_r2 <= din_valid_3_10_r1;

    din_3_10.data <= hash_out_valid_filter_3_10 ? hash_out_3_10 : 0;
    din_3_10.last <= out_new_pkt;
    din_3_10.bucket <= 3;


    din_3_10_r1 <= din_3_10;
    din_3_10_r2 <= din_3_10_r1;
    din_valid_3_11 <= out_new_pkt | hash_out_valid_filter_3_11;
    din_valid_3_11_r1 <= din_valid_3_11;
    din_valid_3_11_r2 <= din_valid_3_11_r1;

    din_3_11.data <= hash_out_valid_filter_3_11 ? hash_out_3_11 : 0;
    din_3_11.last <= out_new_pkt;
    din_3_11.bucket <= 3;


    din_3_11_r1 <= din_3_11;
    din_3_11_r2 <= din_3_11_r1;
    din_valid_3_12 <= out_new_pkt | hash_out_valid_filter_3_12;
    din_valid_3_12_r1 <= din_valid_3_12;
    din_valid_3_12_r2 <= din_valid_3_12_r1;

    din_3_12.data <= hash_out_valid_filter_3_12 ? hash_out_3_12 : 0;
    din_3_12.last <= out_new_pkt;
    din_3_12.bucket <= 3;


    din_3_12_r1 <= din_3_12;
    din_3_12_r2 <= din_3_12_r1;
    din_valid_3_13 <= out_new_pkt | hash_out_valid_filter_3_13;
    din_valid_3_13_r1 <= din_valid_3_13;
    din_valid_3_13_r2 <= din_valid_3_13_r1;

    din_3_13.data <= hash_out_valid_filter_3_13 ? hash_out_3_13 : 0;
    din_3_13.last <= out_new_pkt;
    din_3_13.bucket <= 3;


    din_3_13_r1 <= din_3_13;
    din_3_13_r2 <= din_3_13_r1;
    din_valid_3_14 <= out_new_pkt | hash_out_valid_filter_3_14;
    din_valid_3_14_r1 <= din_valid_3_14;
    din_valid_3_14_r2 <= din_valid_3_14_r1;

    din_3_14.data <= hash_out_valid_filter_3_14 ? hash_out_3_14 : 0;
    din_3_14.last <= out_new_pkt;
    din_3_14.bucket <= 3;


    din_3_14_r1 <= din_3_14;
    din_3_14_r2 <= din_3_14_r1;
    din_valid_3_15 <= out_new_pkt | hash_out_valid_filter_3_15;
    din_valid_3_15_r1 <= din_valid_3_15;
    din_valid_3_15_r2 <= din_valid_3_15_r1;

    din_3_15.data <= hash_out_valid_filter_3_15 ? hash_out_3_15 : 0;
    din_3_15.last <= out_new_pkt;
    din_3_15.bucket <= 3;


    din_3_15_r1 <= din_3_15;
    din_3_15_r2 <= din_3_15_r1;
    din_valid_3_16 <= out_new_pkt | hash_out_valid_filter_3_16;
    din_valid_3_16_r1 <= din_valid_3_16;
    din_valid_3_16_r2 <= din_valid_3_16_r1;

    din_3_16.data <= hash_out_valid_filter_3_16 ? hash_out_3_16 : 0;
    din_3_16.last <= out_new_pkt;
    din_3_16.bucket <= 3;


    din_3_16_r1 <= din_3_16;
    din_3_16_r2 <= din_3_16_r1;
    din_valid_3_17 <= out_new_pkt | hash_out_valid_filter_3_17;
    din_valid_3_17_r1 <= din_valid_3_17;
    din_valid_3_17_r2 <= din_valid_3_17_r1;

    din_3_17.data <= hash_out_valid_filter_3_17 ? hash_out_3_17 : 0;
    din_3_17.last <= out_new_pkt;
    din_3_17.bucket <= 3;


    din_3_17_r1 <= din_3_17;
    din_3_17_r2 <= din_3_17_r1;
    din_valid_3_18 <= out_new_pkt | hash_out_valid_filter_3_18;
    din_valid_3_18_r1 <= din_valid_3_18;
    din_valid_3_18_r2 <= din_valid_3_18_r1;

    din_3_18.data <= hash_out_valid_filter_3_18 ? hash_out_3_18 : 0;
    din_3_18.last <= out_new_pkt;
    din_3_18.bucket <= 3;


    din_3_18_r1 <= din_3_18;
    din_3_18_r2 <= din_3_18_r1;
    din_valid_3_19 <= out_new_pkt | hash_out_valid_filter_3_19;
    din_valid_3_19_r1 <= din_valid_3_19;
    din_valid_3_19_r2 <= din_valid_3_19_r1;

    din_3_19.data <= hash_out_valid_filter_3_19 ? hash_out_3_19 : 0;
    din_3_19.last <= out_new_pkt;
    din_3_19.bucket <= 3;


    din_3_19_r1 <= din_3_19;
    din_3_19_r2 <= din_3_19_r1;
    din_valid_3_20 <= out_new_pkt | hash_out_valid_filter_3_20;
    din_valid_3_20_r1 <= din_valid_3_20;
    din_valid_3_20_r2 <= din_valid_3_20_r1;

    din_3_20.data <= hash_out_valid_filter_3_20 ? hash_out_3_20 : 0;
    din_3_20.last <= out_new_pkt;
    din_3_20.bucket <= 3;


    din_3_20_r1 <= din_3_20;
    din_3_20_r2 <= din_3_20_r1;
    din_valid_3_21 <= out_new_pkt | hash_out_valid_filter_3_21;
    din_valid_3_21_r1 <= din_valid_3_21;
    din_valid_3_21_r2 <= din_valid_3_21_r1;

    din_3_21.data <= hash_out_valid_filter_3_21 ? hash_out_3_21 : 0;
    din_3_21.last <= out_new_pkt;
    din_3_21.bucket <= 3;


    din_3_21_r1 <= din_3_21;
    din_3_21_r2 <= din_3_21_r1;
    din_valid_3_22 <= out_new_pkt | hash_out_valid_filter_3_22;
    din_valid_3_22_r1 <= din_valid_3_22;
    din_valid_3_22_r2 <= din_valid_3_22_r1;

    din_3_22.data <= hash_out_valid_filter_3_22 ? hash_out_3_22 : 0;
    din_3_22.last <= out_new_pkt;
    din_3_22.bucket <= 3;


    din_3_22_r1 <= din_3_22;
    din_3_22_r2 <= din_3_22_r1;
    din_valid_3_23 <= out_new_pkt | hash_out_valid_filter_3_23;
    din_valid_3_23_r1 <= din_valid_3_23;
    din_valid_3_23_r2 <= din_valid_3_23_r1;

    din_3_23.data <= hash_out_valid_filter_3_23 ? hash_out_3_23 : 0;
    din_3_23.last <= out_new_pkt;
    din_3_23.bucket <= 3;


    din_3_23_r1 <= din_3_23;
    din_3_23_r2 <= din_3_23_r1;
    din_valid_3_24 <= out_new_pkt | hash_out_valid_filter_3_24;
    din_valid_3_24_r1 <= din_valid_3_24;
    din_valid_3_24_r2 <= din_valid_3_24_r1;

    din_3_24.data <= hash_out_valid_filter_3_24 ? hash_out_3_24 : 0;
    din_3_24.last <= out_new_pkt;
    din_3_24.bucket <= 3;


    din_3_24_r1 <= din_3_24;
    din_3_24_r2 <= din_3_24_r1;
    din_valid_3_25 <= out_new_pkt | hash_out_valid_filter_3_25;
    din_valid_3_25_r1 <= din_valid_3_25;
    din_valid_3_25_r2 <= din_valid_3_25_r1;

    din_3_25.data <= hash_out_valid_filter_3_25 ? hash_out_3_25 : 0;
    din_3_25.last <= out_new_pkt;
    din_3_25.bucket <= 3;


    din_3_25_r1 <= din_3_25;
    din_3_25_r2 <= din_3_25_r1;
    din_valid_3_26 <= out_new_pkt | hash_out_valid_filter_3_26;
    din_valid_3_26_r1 <= din_valid_3_26;
    din_valid_3_26_r2 <= din_valid_3_26_r1;

    din_3_26.data <= hash_out_valid_filter_3_26 ? hash_out_3_26 : 0;
    din_3_26.last <= out_new_pkt;
    din_3_26.bucket <= 3;


    din_3_26_r1 <= din_3_26;
    din_3_26_r2 <= din_3_26_r1;
    din_valid_3_27 <= out_new_pkt | hash_out_valid_filter_3_27;
    din_valid_3_27_r1 <= din_valid_3_27;
    din_valid_3_27_r2 <= din_valid_3_27_r1;

    din_3_27.data <= hash_out_valid_filter_3_27 ? hash_out_3_27 : 0;
    din_3_27.last <= out_new_pkt;
    din_3_27.bucket <= 3;


    din_3_27_r1 <= din_3_27;
    din_3_27_r2 <= din_3_27_r1;
    din_valid_3_28 <= out_new_pkt | hash_out_valid_filter_3_28;
    din_valid_3_28_r1 <= din_valid_3_28;
    din_valid_3_28_r2 <= din_valid_3_28_r1;

    din_3_28.data <= hash_out_valid_filter_3_28 ? hash_out_3_28 : 0;
    din_3_28.last <= out_new_pkt;
    din_3_28.bucket <= 3;


    din_3_28_r1 <= din_3_28;
    din_3_28_r2 <= din_3_28_r1;
    din_valid_3_29 <= out_new_pkt | hash_out_valid_filter_3_29;
    din_valid_3_29_r1 <= din_valid_3_29;
    din_valid_3_29_r2 <= din_valid_3_29_r1;

    din_3_29.data <= hash_out_valid_filter_3_29 ? hash_out_3_29 : 0;
    din_3_29.last <= out_new_pkt;
    din_3_29.bucket <= 3;


    din_3_29_r1 <= din_3_29;
    din_3_29_r2 <= din_3_29_r1;
    din_valid_3_30 <= out_new_pkt | hash_out_valid_filter_3_30;
    din_valid_3_30_r1 <= din_valid_3_30;
    din_valid_3_30_r2 <= din_valid_3_30_r1;

    din_3_30.data <= hash_out_valid_filter_3_30 ? hash_out_3_30 : 0;
    din_3_30.last <= out_new_pkt;
    din_3_30.bucket <= 3;


    din_3_30_r1 <= din_3_30;
    din_3_30_r2 <= din_3_30_r1;
    din_valid_3_31 <= out_new_pkt | hash_out_valid_filter_3_31;
    din_valid_3_31_r1 <= din_valid_3_31;
    din_valid_3_31_r2 <= din_valid_3_31_r1;

    din_3_31.data <= hash_out_valid_filter_3_31 ? hash_out_3_31 : 0;
    din_3_31.last <= out_new_pkt;
    din_3_31.bucket <= 3;


    din_3_31_r1 <= din_3_31;
    din_3_31_r2 <= din_3_31_r1;
    din_valid_4_0 <= out_new_pkt | hash_out_valid_filter_4_0;
    din_valid_4_0_r1 <= din_valid_4_0;
    din_valid_4_0_r2 <= din_valid_4_0_r1;

    din_4_0.data <= hash_out_valid_filter_4_0 ? hash_out_4_0 : 0;
    din_4_0.last <= out_new_pkt;
    din_4_0.bucket <= 4;


    din_4_0_r1 <= din_4_0;
    din_4_0_r2 <= din_4_0_r1;
    din_valid_4_1 <= out_new_pkt | hash_out_valid_filter_4_1;
    din_valid_4_1_r1 <= din_valid_4_1;
    din_valid_4_1_r2 <= din_valid_4_1_r1;

    din_4_1.data <= hash_out_valid_filter_4_1 ? hash_out_4_1 : 0;
    din_4_1.last <= out_new_pkt;
    din_4_1.bucket <= 4;


    din_4_1_r1 <= din_4_1;
    din_4_1_r2 <= din_4_1_r1;
    din_valid_4_2 <= out_new_pkt | hash_out_valid_filter_4_2;
    din_valid_4_2_r1 <= din_valid_4_2;
    din_valid_4_2_r2 <= din_valid_4_2_r1;

    din_4_2.data <= hash_out_valid_filter_4_2 ? hash_out_4_2 : 0;
    din_4_2.last <= out_new_pkt;
    din_4_2.bucket <= 4;


    din_4_2_r1 <= din_4_2;
    din_4_2_r2 <= din_4_2_r1;
    din_valid_4_3 <= out_new_pkt | hash_out_valid_filter_4_3;
    din_valid_4_3_r1 <= din_valid_4_3;
    din_valid_4_3_r2 <= din_valid_4_3_r1;

    din_4_3.data <= hash_out_valid_filter_4_3 ? hash_out_4_3 : 0;
    din_4_3.last <= out_new_pkt;
    din_4_3.bucket <= 4;


    din_4_3_r1 <= din_4_3;
    din_4_3_r2 <= din_4_3_r1;
    din_valid_4_4 <= out_new_pkt | hash_out_valid_filter_4_4;
    din_valid_4_4_r1 <= din_valid_4_4;
    din_valid_4_4_r2 <= din_valid_4_4_r1;

    din_4_4.data <= hash_out_valid_filter_4_4 ? hash_out_4_4 : 0;
    din_4_4.last <= out_new_pkt;
    din_4_4.bucket <= 4;


    din_4_4_r1 <= din_4_4;
    din_4_4_r2 <= din_4_4_r1;
    din_valid_4_5 <= out_new_pkt | hash_out_valid_filter_4_5;
    din_valid_4_5_r1 <= din_valid_4_5;
    din_valid_4_5_r2 <= din_valid_4_5_r1;

    din_4_5.data <= hash_out_valid_filter_4_5 ? hash_out_4_5 : 0;
    din_4_5.last <= out_new_pkt;
    din_4_5.bucket <= 4;


    din_4_5_r1 <= din_4_5;
    din_4_5_r2 <= din_4_5_r1;
    din_valid_4_6 <= out_new_pkt | hash_out_valid_filter_4_6;
    din_valid_4_6_r1 <= din_valid_4_6;
    din_valid_4_6_r2 <= din_valid_4_6_r1;

    din_4_6.data <= hash_out_valid_filter_4_6 ? hash_out_4_6 : 0;
    din_4_6.last <= out_new_pkt;
    din_4_6.bucket <= 4;


    din_4_6_r1 <= din_4_6;
    din_4_6_r2 <= din_4_6_r1;
    din_valid_4_7 <= out_new_pkt | hash_out_valid_filter_4_7;
    din_valid_4_7_r1 <= din_valid_4_7;
    din_valid_4_7_r2 <= din_valid_4_7_r1;

    din_4_7.data <= hash_out_valid_filter_4_7 ? hash_out_4_7 : 0;
    din_4_7.last <= out_new_pkt;
    din_4_7.bucket <= 4;


    din_4_7_r1 <= din_4_7;
    din_4_7_r2 <= din_4_7_r1;
    din_valid_4_8 <= out_new_pkt | hash_out_valid_filter_4_8;
    din_valid_4_8_r1 <= din_valid_4_8;
    din_valid_4_8_r2 <= din_valid_4_8_r1;

    din_4_8.data <= hash_out_valid_filter_4_8 ? hash_out_4_8 : 0;
    din_4_8.last <= out_new_pkt;
    din_4_8.bucket <= 4;


    din_4_8_r1 <= din_4_8;
    din_4_8_r2 <= din_4_8_r1;
    din_valid_4_9 <= out_new_pkt | hash_out_valid_filter_4_9;
    din_valid_4_9_r1 <= din_valid_4_9;
    din_valid_4_9_r2 <= din_valid_4_9_r1;

    din_4_9.data <= hash_out_valid_filter_4_9 ? hash_out_4_9 : 0;
    din_4_9.last <= out_new_pkt;
    din_4_9.bucket <= 4;


    din_4_9_r1 <= din_4_9;
    din_4_9_r2 <= din_4_9_r1;
    din_valid_4_10 <= out_new_pkt | hash_out_valid_filter_4_10;
    din_valid_4_10_r1 <= din_valid_4_10;
    din_valid_4_10_r2 <= din_valid_4_10_r1;

    din_4_10.data <= hash_out_valid_filter_4_10 ? hash_out_4_10 : 0;
    din_4_10.last <= out_new_pkt;
    din_4_10.bucket <= 4;


    din_4_10_r1 <= din_4_10;
    din_4_10_r2 <= din_4_10_r1;
    din_valid_4_11 <= out_new_pkt | hash_out_valid_filter_4_11;
    din_valid_4_11_r1 <= din_valid_4_11;
    din_valid_4_11_r2 <= din_valid_4_11_r1;

    din_4_11.data <= hash_out_valid_filter_4_11 ? hash_out_4_11 : 0;
    din_4_11.last <= out_new_pkt;
    din_4_11.bucket <= 4;


    din_4_11_r1 <= din_4_11;
    din_4_11_r2 <= din_4_11_r1;
    din_valid_4_12 <= out_new_pkt | hash_out_valid_filter_4_12;
    din_valid_4_12_r1 <= din_valid_4_12;
    din_valid_4_12_r2 <= din_valid_4_12_r1;

    din_4_12.data <= hash_out_valid_filter_4_12 ? hash_out_4_12 : 0;
    din_4_12.last <= out_new_pkt;
    din_4_12.bucket <= 4;


    din_4_12_r1 <= din_4_12;
    din_4_12_r2 <= din_4_12_r1;
    din_valid_4_13 <= out_new_pkt | hash_out_valid_filter_4_13;
    din_valid_4_13_r1 <= din_valid_4_13;
    din_valid_4_13_r2 <= din_valid_4_13_r1;

    din_4_13.data <= hash_out_valid_filter_4_13 ? hash_out_4_13 : 0;
    din_4_13.last <= out_new_pkt;
    din_4_13.bucket <= 4;


    din_4_13_r1 <= din_4_13;
    din_4_13_r2 <= din_4_13_r1;
    din_valid_4_14 <= out_new_pkt | hash_out_valid_filter_4_14;
    din_valid_4_14_r1 <= din_valid_4_14;
    din_valid_4_14_r2 <= din_valid_4_14_r1;

    din_4_14.data <= hash_out_valid_filter_4_14 ? hash_out_4_14 : 0;
    din_4_14.last <= out_new_pkt;
    din_4_14.bucket <= 4;


    din_4_14_r1 <= din_4_14;
    din_4_14_r2 <= din_4_14_r1;
    din_valid_4_15 <= out_new_pkt | hash_out_valid_filter_4_15;
    din_valid_4_15_r1 <= din_valid_4_15;
    din_valid_4_15_r2 <= din_valid_4_15_r1;

    din_4_15.data <= hash_out_valid_filter_4_15 ? hash_out_4_15 : 0;
    din_4_15.last <= out_new_pkt;
    din_4_15.bucket <= 4;


    din_4_15_r1 <= din_4_15;
    din_4_15_r2 <= din_4_15_r1;
    din_valid_4_16 <= out_new_pkt | hash_out_valid_filter_4_16;
    din_valid_4_16_r1 <= din_valid_4_16;
    din_valid_4_16_r2 <= din_valid_4_16_r1;

    din_4_16.data <= hash_out_valid_filter_4_16 ? hash_out_4_16 : 0;
    din_4_16.last <= out_new_pkt;
    din_4_16.bucket <= 4;


    din_4_16_r1 <= din_4_16;
    din_4_16_r2 <= din_4_16_r1;
    din_valid_4_17 <= out_new_pkt | hash_out_valid_filter_4_17;
    din_valid_4_17_r1 <= din_valid_4_17;
    din_valid_4_17_r2 <= din_valid_4_17_r1;

    din_4_17.data <= hash_out_valid_filter_4_17 ? hash_out_4_17 : 0;
    din_4_17.last <= out_new_pkt;
    din_4_17.bucket <= 4;


    din_4_17_r1 <= din_4_17;
    din_4_17_r2 <= din_4_17_r1;
    din_valid_4_18 <= out_new_pkt | hash_out_valid_filter_4_18;
    din_valid_4_18_r1 <= din_valid_4_18;
    din_valid_4_18_r2 <= din_valid_4_18_r1;

    din_4_18.data <= hash_out_valid_filter_4_18 ? hash_out_4_18 : 0;
    din_4_18.last <= out_new_pkt;
    din_4_18.bucket <= 4;


    din_4_18_r1 <= din_4_18;
    din_4_18_r2 <= din_4_18_r1;
    din_valid_4_19 <= out_new_pkt | hash_out_valid_filter_4_19;
    din_valid_4_19_r1 <= din_valid_4_19;
    din_valid_4_19_r2 <= din_valid_4_19_r1;

    din_4_19.data <= hash_out_valid_filter_4_19 ? hash_out_4_19 : 0;
    din_4_19.last <= out_new_pkt;
    din_4_19.bucket <= 4;


    din_4_19_r1 <= din_4_19;
    din_4_19_r2 <= din_4_19_r1;
    din_valid_4_20 <= out_new_pkt | hash_out_valid_filter_4_20;
    din_valid_4_20_r1 <= din_valid_4_20;
    din_valid_4_20_r2 <= din_valid_4_20_r1;

    din_4_20.data <= hash_out_valid_filter_4_20 ? hash_out_4_20 : 0;
    din_4_20.last <= out_new_pkt;
    din_4_20.bucket <= 4;


    din_4_20_r1 <= din_4_20;
    din_4_20_r2 <= din_4_20_r1;
    din_valid_4_21 <= out_new_pkt | hash_out_valid_filter_4_21;
    din_valid_4_21_r1 <= din_valid_4_21;
    din_valid_4_21_r2 <= din_valid_4_21_r1;

    din_4_21.data <= hash_out_valid_filter_4_21 ? hash_out_4_21 : 0;
    din_4_21.last <= out_new_pkt;
    din_4_21.bucket <= 4;


    din_4_21_r1 <= din_4_21;
    din_4_21_r2 <= din_4_21_r1;
    din_valid_4_22 <= out_new_pkt | hash_out_valid_filter_4_22;
    din_valid_4_22_r1 <= din_valid_4_22;
    din_valid_4_22_r2 <= din_valid_4_22_r1;

    din_4_22.data <= hash_out_valid_filter_4_22 ? hash_out_4_22 : 0;
    din_4_22.last <= out_new_pkt;
    din_4_22.bucket <= 4;


    din_4_22_r1 <= din_4_22;
    din_4_22_r2 <= din_4_22_r1;
    din_valid_4_23 <= out_new_pkt | hash_out_valid_filter_4_23;
    din_valid_4_23_r1 <= din_valid_4_23;
    din_valid_4_23_r2 <= din_valid_4_23_r1;

    din_4_23.data <= hash_out_valid_filter_4_23 ? hash_out_4_23 : 0;
    din_4_23.last <= out_new_pkt;
    din_4_23.bucket <= 4;


    din_4_23_r1 <= din_4_23;
    din_4_23_r2 <= din_4_23_r1;
    din_valid_4_24 <= out_new_pkt | hash_out_valid_filter_4_24;
    din_valid_4_24_r1 <= din_valid_4_24;
    din_valid_4_24_r2 <= din_valid_4_24_r1;

    din_4_24.data <= hash_out_valid_filter_4_24 ? hash_out_4_24 : 0;
    din_4_24.last <= out_new_pkt;
    din_4_24.bucket <= 4;


    din_4_24_r1 <= din_4_24;
    din_4_24_r2 <= din_4_24_r1;
    din_valid_4_25 <= out_new_pkt | hash_out_valid_filter_4_25;
    din_valid_4_25_r1 <= din_valid_4_25;
    din_valid_4_25_r2 <= din_valid_4_25_r1;

    din_4_25.data <= hash_out_valid_filter_4_25 ? hash_out_4_25 : 0;
    din_4_25.last <= out_new_pkt;
    din_4_25.bucket <= 4;


    din_4_25_r1 <= din_4_25;
    din_4_25_r2 <= din_4_25_r1;
    din_valid_4_26 <= out_new_pkt | hash_out_valid_filter_4_26;
    din_valid_4_26_r1 <= din_valid_4_26;
    din_valid_4_26_r2 <= din_valid_4_26_r1;

    din_4_26.data <= hash_out_valid_filter_4_26 ? hash_out_4_26 : 0;
    din_4_26.last <= out_new_pkt;
    din_4_26.bucket <= 4;


    din_4_26_r1 <= din_4_26;
    din_4_26_r2 <= din_4_26_r1;
    din_valid_4_27 <= out_new_pkt | hash_out_valid_filter_4_27;
    din_valid_4_27_r1 <= din_valid_4_27;
    din_valid_4_27_r2 <= din_valid_4_27_r1;

    din_4_27.data <= hash_out_valid_filter_4_27 ? hash_out_4_27 : 0;
    din_4_27.last <= out_new_pkt;
    din_4_27.bucket <= 4;


    din_4_27_r1 <= din_4_27;
    din_4_27_r2 <= din_4_27_r1;
    din_valid_4_28 <= out_new_pkt | hash_out_valid_filter_4_28;
    din_valid_4_28_r1 <= din_valid_4_28;
    din_valid_4_28_r2 <= din_valid_4_28_r1;

    din_4_28.data <= hash_out_valid_filter_4_28 ? hash_out_4_28 : 0;
    din_4_28.last <= out_new_pkt;
    din_4_28.bucket <= 4;


    din_4_28_r1 <= din_4_28;
    din_4_28_r2 <= din_4_28_r1;
    din_valid_4_29 <= out_new_pkt | hash_out_valid_filter_4_29;
    din_valid_4_29_r1 <= din_valid_4_29;
    din_valid_4_29_r2 <= din_valid_4_29_r1;

    din_4_29.data <= hash_out_valid_filter_4_29 ? hash_out_4_29 : 0;
    din_4_29.last <= out_new_pkt;
    din_4_29.bucket <= 4;


    din_4_29_r1 <= din_4_29;
    din_4_29_r2 <= din_4_29_r1;
    din_valid_4_30 <= out_new_pkt | hash_out_valid_filter_4_30;
    din_valid_4_30_r1 <= din_valid_4_30;
    din_valid_4_30_r2 <= din_valid_4_30_r1;

    din_4_30.data <= hash_out_valid_filter_4_30 ? hash_out_4_30 : 0;
    din_4_30.last <= out_new_pkt;
    din_4_30.bucket <= 4;


    din_4_30_r1 <= din_4_30;
    din_4_30_r2 <= din_4_30_r1;
    din_valid_4_31 <= out_new_pkt | hash_out_valid_filter_4_31;
    din_valid_4_31_r1 <= din_valid_4_31;
    din_valid_4_31_r2 <= din_valid_4_31_r1;

    din_4_31.data <= hash_out_valid_filter_4_31 ? hash_out_4_31 : 0;
    din_4_31.last <= out_new_pkt;
    din_4_31.bucket <= 4;


    din_4_31_r1 <= din_4_31;
    din_4_31_r2 <= din_4_31_r1;
    din_valid_5_0 <= out_new_pkt | hash_out_valid_filter_5_0;
    din_valid_5_0_r1 <= din_valid_5_0;
    din_valid_5_0_r2 <= din_valid_5_0_r1;

    din_5_0.data <= hash_out_valid_filter_5_0 ? hash_out_5_0 : 0;
    din_5_0.last <= out_new_pkt;
    din_5_0.bucket <= 5;


    din_5_0_r1 <= din_5_0;
    din_5_0_r2 <= din_5_0_r1;
    din_valid_5_1 <= out_new_pkt | hash_out_valid_filter_5_1;
    din_valid_5_1_r1 <= din_valid_5_1;
    din_valid_5_1_r2 <= din_valid_5_1_r1;

    din_5_1.data <= hash_out_valid_filter_5_1 ? hash_out_5_1 : 0;
    din_5_1.last <= out_new_pkt;
    din_5_1.bucket <= 5;


    din_5_1_r1 <= din_5_1;
    din_5_1_r2 <= din_5_1_r1;
    din_valid_5_2 <= out_new_pkt | hash_out_valid_filter_5_2;
    din_valid_5_2_r1 <= din_valid_5_2;
    din_valid_5_2_r2 <= din_valid_5_2_r1;

    din_5_2.data <= hash_out_valid_filter_5_2 ? hash_out_5_2 : 0;
    din_5_2.last <= out_new_pkt;
    din_5_2.bucket <= 5;


    din_5_2_r1 <= din_5_2;
    din_5_2_r2 <= din_5_2_r1;
    din_valid_5_3 <= out_new_pkt | hash_out_valid_filter_5_3;
    din_valid_5_3_r1 <= din_valid_5_3;
    din_valid_5_3_r2 <= din_valid_5_3_r1;

    din_5_3.data <= hash_out_valid_filter_5_3 ? hash_out_5_3 : 0;
    din_5_3.last <= out_new_pkt;
    din_5_3.bucket <= 5;


    din_5_3_r1 <= din_5_3;
    din_5_3_r2 <= din_5_3_r1;
    din_valid_5_4 <= out_new_pkt | hash_out_valid_filter_5_4;
    din_valid_5_4_r1 <= din_valid_5_4;
    din_valid_5_4_r2 <= din_valid_5_4_r1;

    din_5_4.data <= hash_out_valid_filter_5_4 ? hash_out_5_4 : 0;
    din_5_4.last <= out_new_pkt;
    din_5_4.bucket <= 5;


    din_5_4_r1 <= din_5_4;
    din_5_4_r2 <= din_5_4_r1;
    din_valid_5_5 <= out_new_pkt | hash_out_valid_filter_5_5;
    din_valid_5_5_r1 <= din_valid_5_5;
    din_valid_5_5_r2 <= din_valid_5_5_r1;

    din_5_5.data <= hash_out_valid_filter_5_5 ? hash_out_5_5 : 0;
    din_5_5.last <= out_new_pkt;
    din_5_5.bucket <= 5;


    din_5_5_r1 <= din_5_5;
    din_5_5_r2 <= din_5_5_r1;
    din_valid_5_6 <= out_new_pkt | hash_out_valid_filter_5_6;
    din_valid_5_6_r1 <= din_valid_5_6;
    din_valid_5_6_r2 <= din_valid_5_6_r1;

    din_5_6.data <= hash_out_valid_filter_5_6 ? hash_out_5_6 : 0;
    din_5_6.last <= out_new_pkt;
    din_5_6.bucket <= 5;


    din_5_6_r1 <= din_5_6;
    din_5_6_r2 <= din_5_6_r1;
    din_valid_5_7 <= out_new_pkt | hash_out_valid_filter_5_7;
    din_valid_5_7_r1 <= din_valid_5_7;
    din_valid_5_7_r2 <= din_valid_5_7_r1;

    din_5_7.data <= hash_out_valid_filter_5_7 ? hash_out_5_7 : 0;
    din_5_7.last <= out_new_pkt;
    din_5_7.bucket <= 5;


    din_5_7_r1 <= din_5_7;
    din_5_7_r2 <= din_5_7_r1;
    din_valid_5_8 <= out_new_pkt | hash_out_valid_filter_5_8;
    din_valid_5_8_r1 <= din_valid_5_8;
    din_valid_5_8_r2 <= din_valid_5_8_r1;

    din_5_8.data <= hash_out_valid_filter_5_8 ? hash_out_5_8 : 0;
    din_5_8.last <= out_new_pkt;
    din_5_8.bucket <= 5;


    din_5_8_r1 <= din_5_8;
    din_5_8_r2 <= din_5_8_r1;
    din_valid_5_9 <= out_new_pkt | hash_out_valid_filter_5_9;
    din_valid_5_9_r1 <= din_valid_5_9;
    din_valid_5_9_r2 <= din_valid_5_9_r1;

    din_5_9.data <= hash_out_valid_filter_5_9 ? hash_out_5_9 : 0;
    din_5_9.last <= out_new_pkt;
    din_5_9.bucket <= 5;


    din_5_9_r1 <= din_5_9;
    din_5_9_r2 <= din_5_9_r1;
    din_valid_5_10 <= out_new_pkt | hash_out_valid_filter_5_10;
    din_valid_5_10_r1 <= din_valid_5_10;
    din_valid_5_10_r2 <= din_valid_5_10_r1;

    din_5_10.data <= hash_out_valid_filter_5_10 ? hash_out_5_10 : 0;
    din_5_10.last <= out_new_pkt;
    din_5_10.bucket <= 5;


    din_5_10_r1 <= din_5_10;
    din_5_10_r2 <= din_5_10_r1;
    din_valid_5_11 <= out_new_pkt | hash_out_valid_filter_5_11;
    din_valid_5_11_r1 <= din_valid_5_11;
    din_valid_5_11_r2 <= din_valid_5_11_r1;

    din_5_11.data <= hash_out_valid_filter_5_11 ? hash_out_5_11 : 0;
    din_5_11.last <= out_new_pkt;
    din_5_11.bucket <= 5;


    din_5_11_r1 <= din_5_11;
    din_5_11_r2 <= din_5_11_r1;
    din_valid_5_12 <= out_new_pkt | hash_out_valid_filter_5_12;
    din_valid_5_12_r1 <= din_valid_5_12;
    din_valid_5_12_r2 <= din_valid_5_12_r1;

    din_5_12.data <= hash_out_valid_filter_5_12 ? hash_out_5_12 : 0;
    din_5_12.last <= out_new_pkt;
    din_5_12.bucket <= 5;


    din_5_12_r1 <= din_5_12;
    din_5_12_r2 <= din_5_12_r1;
    din_valid_5_13 <= out_new_pkt | hash_out_valid_filter_5_13;
    din_valid_5_13_r1 <= din_valid_5_13;
    din_valid_5_13_r2 <= din_valid_5_13_r1;

    din_5_13.data <= hash_out_valid_filter_5_13 ? hash_out_5_13 : 0;
    din_5_13.last <= out_new_pkt;
    din_5_13.bucket <= 5;


    din_5_13_r1 <= din_5_13;
    din_5_13_r2 <= din_5_13_r1;
    din_valid_5_14 <= out_new_pkt | hash_out_valid_filter_5_14;
    din_valid_5_14_r1 <= din_valid_5_14;
    din_valid_5_14_r2 <= din_valid_5_14_r1;

    din_5_14.data <= hash_out_valid_filter_5_14 ? hash_out_5_14 : 0;
    din_5_14.last <= out_new_pkt;
    din_5_14.bucket <= 5;


    din_5_14_r1 <= din_5_14;
    din_5_14_r2 <= din_5_14_r1;
    din_valid_5_15 <= out_new_pkt | hash_out_valid_filter_5_15;
    din_valid_5_15_r1 <= din_valid_5_15;
    din_valid_5_15_r2 <= din_valid_5_15_r1;

    din_5_15.data <= hash_out_valid_filter_5_15 ? hash_out_5_15 : 0;
    din_5_15.last <= out_new_pkt;
    din_5_15.bucket <= 5;


    din_5_15_r1 <= din_5_15;
    din_5_15_r2 <= din_5_15_r1;
    din_valid_5_16 <= out_new_pkt | hash_out_valid_filter_5_16;
    din_valid_5_16_r1 <= din_valid_5_16;
    din_valid_5_16_r2 <= din_valid_5_16_r1;

    din_5_16.data <= hash_out_valid_filter_5_16 ? hash_out_5_16 : 0;
    din_5_16.last <= out_new_pkt;
    din_5_16.bucket <= 5;


    din_5_16_r1 <= din_5_16;
    din_5_16_r2 <= din_5_16_r1;
    din_valid_5_17 <= out_new_pkt | hash_out_valid_filter_5_17;
    din_valid_5_17_r1 <= din_valid_5_17;
    din_valid_5_17_r2 <= din_valid_5_17_r1;

    din_5_17.data <= hash_out_valid_filter_5_17 ? hash_out_5_17 : 0;
    din_5_17.last <= out_new_pkt;
    din_5_17.bucket <= 5;


    din_5_17_r1 <= din_5_17;
    din_5_17_r2 <= din_5_17_r1;
    din_valid_5_18 <= out_new_pkt | hash_out_valid_filter_5_18;
    din_valid_5_18_r1 <= din_valid_5_18;
    din_valid_5_18_r2 <= din_valid_5_18_r1;

    din_5_18.data <= hash_out_valid_filter_5_18 ? hash_out_5_18 : 0;
    din_5_18.last <= out_new_pkt;
    din_5_18.bucket <= 5;


    din_5_18_r1 <= din_5_18;
    din_5_18_r2 <= din_5_18_r1;
    din_valid_5_19 <= out_new_pkt | hash_out_valid_filter_5_19;
    din_valid_5_19_r1 <= din_valid_5_19;
    din_valid_5_19_r2 <= din_valid_5_19_r1;

    din_5_19.data <= hash_out_valid_filter_5_19 ? hash_out_5_19 : 0;
    din_5_19.last <= out_new_pkt;
    din_5_19.bucket <= 5;


    din_5_19_r1 <= din_5_19;
    din_5_19_r2 <= din_5_19_r1;
    din_valid_5_20 <= out_new_pkt | hash_out_valid_filter_5_20;
    din_valid_5_20_r1 <= din_valid_5_20;
    din_valid_5_20_r2 <= din_valid_5_20_r1;

    din_5_20.data <= hash_out_valid_filter_5_20 ? hash_out_5_20 : 0;
    din_5_20.last <= out_new_pkt;
    din_5_20.bucket <= 5;


    din_5_20_r1 <= din_5_20;
    din_5_20_r2 <= din_5_20_r1;
    din_valid_5_21 <= out_new_pkt | hash_out_valid_filter_5_21;
    din_valid_5_21_r1 <= din_valid_5_21;
    din_valid_5_21_r2 <= din_valid_5_21_r1;

    din_5_21.data <= hash_out_valid_filter_5_21 ? hash_out_5_21 : 0;
    din_5_21.last <= out_new_pkt;
    din_5_21.bucket <= 5;


    din_5_21_r1 <= din_5_21;
    din_5_21_r2 <= din_5_21_r1;
    din_valid_5_22 <= out_new_pkt | hash_out_valid_filter_5_22;
    din_valid_5_22_r1 <= din_valid_5_22;
    din_valid_5_22_r2 <= din_valid_5_22_r1;

    din_5_22.data <= hash_out_valid_filter_5_22 ? hash_out_5_22 : 0;
    din_5_22.last <= out_new_pkt;
    din_5_22.bucket <= 5;


    din_5_22_r1 <= din_5_22;
    din_5_22_r2 <= din_5_22_r1;
    din_valid_5_23 <= out_new_pkt | hash_out_valid_filter_5_23;
    din_valid_5_23_r1 <= din_valid_5_23;
    din_valid_5_23_r2 <= din_valid_5_23_r1;

    din_5_23.data <= hash_out_valid_filter_5_23 ? hash_out_5_23 : 0;
    din_5_23.last <= out_new_pkt;
    din_5_23.bucket <= 5;


    din_5_23_r1 <= din_5_23;
    din_5_23_r2 <= din_5_23_r1;
    din_valid_5_24 <= out_new_pkt | hash_out_valid_filter_5_24;
    din_valid_5_24_r1 <= din_valid_5_24;
    din_valid_5_24_r2 <= din_valid_5_24_r1;

    din_5_24.data <= hash_out_valid_filter_5_24 ? hash_out_5_24 : 0;
    din_5_24.last <= out_new_pkt;
    din_5_24.bucket <= 5;


    din_5_24_r1 <= din_5_24;
    din_5_24_r2 <= din_5_24_r1;
    din_valid_5_25 <= out_new_pkt | hash_out_valid_filter_5_25;
    din_valid_5_25_r1 <= din_valid_5_25;
    din_valid_5_25_r2 <= din_valid_5_25_r1;

    din_5_25.data <= hash_out_valid_filter_5_25 ? hash_out_5_25 : 0;
    din_5_25.last <= out_new_pkt;
    din_5_25.bucket <= 5;


    din_5_25_r1 <= din_5_25;
    din_5_25_r2 <= din_5_25_r1;
    din_valid_5_26 <= out_new_pkt | hash_out_valid_filter_5_26;
    din_valid_5_26_r1 <= din_valid_5_26;
    din_valid_5_26_r2 <= din_valid_5_26_r1;

    din_5_26.data <= hash_out_valid_filter_5_26 ? hash_out_5_26 : 0;
    din_5_26.last <= out_new_pkt;
    din_5_26.bucket <= 5;


    din_5_26_r1 <= din_5_26;
    din_5_26_r2 <= din_5_26_r1;
    din_valid_5_27 <= out_new_pkt | hash_out_valid_filter_5_27;
    din_valid_5_27_r1 <= din_valid_5_27;
    din_valid_5_27_r2 <= din_valid_5_27_r1;

    din_5_27.data <= hash_out_valid_filter_5_27 ? hash_out_5_27 : 0;
    din_5_27.last <= out_new_pkt;
    din_5_27.bucket <= 5;


    din_5_27_r1 <= din_5_27;
    din_5_27_r2 <= din_5_27_r1;
    din_valid_5_28 <= out_new_pkt | hash_out_valid_filter_5_28;
    din_valid_5_28_r1 <= din_valid_5_28;
    din_valid_5_28_r2 <= din_valid_5_28_r1;

    din_5_28.data <= hash_out_valid_filter_5_28 ? hash_out_5_28 : 0;
    din_5_28.last <= out_new_pkt;
    din_5_28.bucket <= 5;


    din_5_28_r1 <= din_5_28;
    din_5_28_r2 <= din_5_28_r1;
    din_valid_5_29 <= out_new_pkt | hash_out_valid_filter_5_29;
    din_valid_5_29_r1 <= din_valid_5_29;
    din_valid_5_29_r2 <= din_valid_5_29_r1;

    din_5_29.data <= hash_out_valid_filter_5_29 ? hash_out_5_29 : 0;
    din_5_29.last <= out_new_pkt;
    din_5_29.bucket <= 5;


    din_5_29_r1 <= din_5_29;
    din_5_29_r2 <= din_5_29_r1;
    din_valid_5_30 <= out_new_pkt | hash_out_valid_filter_5_30;
    din_valid_5_30_r1 <= din_valid_5_30;
    din_valid_5_30_r2 <= din_valid_5_30_r1;

    din_5_30.data <= hash_out_valid_filter_5_30 ? hash_out_5_30 : 0;
    din_5_30.last <= out_new_pkt;
    din_5_30.bucket <= 5;


    din_5_30_r1 <= din_5_30;
    din_5_30_r2 <= din_5_30_r1;
    din_valid_5_31 <= out_new_pkt | hash_out_valid_filter_5_31;
    din_valid_5_31_r1 <= din_valid_5_31;
    din_valid_5_31_r2 <= din_valid_5_31_r1;

    din_5_31.data <= hash_out_valid_filter_5_31 ? hash_out_5_31 : 0;
    din_5_31.last <= out_new_pkt;
    din_5_31.bucket <= 5;


    din_5_31_r1 <= din_5_31;
    din_5_31_r2 <= din_5_31_r1;
    din_valid_6_0 <= out_new_pkt | hash_out_valid_filter_6_0;
    din_valid_6_0_r1 <= din_valid_6_0;
    din_valid_6_0_r2 <= din_valid_6_0_r1;

    din_6_0.data <= hash_out_valid_filter_6_0 ? hash_out_6_0 : 0;
    din_6_0.last <= out_new_pkt;
    din_6_0.bucket <= 6;


    din_6_0_r1 <= din_6_0;
    din_6_0_r2 <= din_6_0_r1;
    din_valid_6_1 <= out_new_pkt | hash_out_valid_filter_6_1;
    din_valid_6_1_r1 <= din_valid_6_1;
    din_valid_6_1_r2 <= din_valid_6_1_r1;

    din_6_1.data <= hash_out_valid_filter_6_1 ? hash_out_6_1 : 0;
    din_6_1.last <= out_new_pkt;
    din_6_1.bucket <= 6;


    din_6_1_r1 <= din_6_1;
    din_6_1_r2 <= din_6_1_r1;
    din_valid_6_2 <= out_new_pkt | hash_out_valid_filter_6_2;
    din_valid_6_2_r1 <= din_valid_6_2;
    din_valid_6_2_r2 <= din_valid_6_2_r1;

    din_6_2.data <= hash_out_valid_filter_6_2 ? hash_out_6_2 : 0;
    din_6_2.last <= out_new_pkt;
    din_6_2.bucket <= 6;


    din_6_2_r1 <= din_6_2;
    din_6_2_r2 <= din_6_2_r1;
    din_valid_6_3 <= out_new_pkt | hash_out_valid_filter_6_3;
    din_valid_6_3_r1 <= din_valid_6_3;
    din_valid_6_3_r2 <= din_valid_6_3_r1;

    din_6_3.data <= hash_out_valid_filter_6_3 ? hash_out_6_3 : 0;
    din_6_3.last <= out_new_pkt;
    din_6_3.bucket <= 6;


    din_6_3_r1 <= din_6_3;
    din_6_3_r2 <= din_6_3_r1;
    din_valid_6_4 <= out_new_pkt | hash_out_valid_filter_6_4;
    din_valid_6_4_r1 <= din_valid_6_4;
    din_valid_6_4_r2 <= din_valid_6_4_r1;

    din_6_4.data <= hash_out_valid_filter_6_4 ? hash_out_6_4 : 0;
    din_6_4.last <= out_new_pkt;
    din_6_4.bucket <= 6;


    din_6_4_r1 <= din_6_4;
    din_6_4_r2 <= din_6_4_r1;
    din_valid_6_5 <= out_new_pkt | hash_out_valid_filter_6_5;
    din_valid_6_5_r1 <= din_valid_6_5;
    din_valid_6_5_r2 <= din_valid_6_5_r1;

    din_6_5.data <= hash_out_valid_filter_6_5 ? hash_out_6_5 : 0;
    din_6_5.last <= out_new_pkt;
    din_6_5.bucket <= 6;


    din_6_5_r1 <= din_6_5;
    din_6_5_r2 <= din_6_5_r1;
    din_valid_6_6 <= out_new_pkt | hash_out_valid_filter_6_6;
    din_valid_6_6_r1 <= din_valid_6_6;
    din_valid_6_6_r2 <= din_valid_6_6_r1;

    din_6_6.data <= hash_out_valid_filter_6_6 ? hash_out_6_6 : 0;
    din_6_6.last <= out_new_pkt;
    din_6_6.bucket <= 6;


    din_6_6_r1 <= din_6_6;
    din_6_6_r2 <= din_6_6_r1;
    din_valid_6_7 <= out_new_pkt | hash_out_valid_filter_6_7;
    din_valid_6_7_r1 <= din_valid_6_7;
    din_valid_6_7_r2 <= din_valid_6_7_r1;

    din_6_7.data <= hash_out_valid_filter_6_7 ? hash_out_6_7 : 0;
    din_6_7.last <= out_new_pkt;
    din_6_7.bucket <= 6;


    din_6_7_r1 <= din_6_7;
    din_6_7_r2 <= din_6_7_r1;
    din_valid_6_8 <= out_new_pkt | hash_out_valid_filter_6_8;
    din_valid_6_8_r1 <= din_valid_6_8;
    din_valid_6_8_r2 <= din_valid_6_8_r1;

    din_6_8.data <= hash_out_valid_filter_6_8 ? hash_out_6_8 : 0;
    din_6_8.last <= out_new_pkt;
    din_6_8.bucket <= 6;


    din_6_8_r1 <= din_6_8;
    din_6_8_r2 <= din_6_8_r1;
    din_valid_6_9 <= out_new_pkt | hash_out_valid_filter_6_9;
    din_valid_6_9_r1 <= din_valid_6_9;
    din_valid_6_9_r2 <= din_valid_6_9_r1;

    din_6_9.data <= hash_out_valid_filter_6_9 ? hash_out_6_9 : 0;
    din_6_9.last <= out_new_pkt;
    din_6_9.bucket <= 6;


    din_6_9_r1 <= din_6_9;
    din_6_9_r2 <= din_6_9_r1;
    din_valid_6_10 <= out_new_pkt | hash_out_valid_filter_6_10;
    din_valid_6_10_r1 <= din_valid_6_10;
    din_valid_6_10_r2 <= din_valid_6_10_r1;

    din_6_10.data <= hash_out_valid_filter_6_10 ? hash_out_6_10 : 0;
    din_6_10.last <= out_new_pkt;
    din_6_10.bucket <= 6;


    din_6_10_r1 <= din_6_10;
    din_6_10_r2 <= din_6_10_r1;
    din_valid_6_11 <= out_new_pkt | hash_out_valid_filter_6_11;
    din_valid_6_11_r1 <= din_valid_6_11;
    din_valid_6_11_r2 <= din_valid_6_11_r1;

    din_6_11.data <= hash_out_valid_filter_6_11 ? hash_out_6_11 : 0;
    din_6_11.last <= out_new_pkt;
    din_6_11.bucket <= 6;


    din_6_11_r1 <= din_6_11;
    din_6_11_r2 <= din_6_11_r1;
    din_valid_6_12 <= out_new_pkt | hash_out_valid_filter_6_12;
    din_valid_6_12_r1 <= din_valid_6_12;
    din_valid_6_12_r2 <= din_valid_6_12_r1;

    din_6_12.data <= hash_out_valid_filter_6_12 ? hash_out_6_12 : 0;
    din_6_12.last <= out_new_pkt;
    din_6_12.bucket <= 6;


    din_6_12_r1 <= din_6_12;
    din_6_12_r2 <= din_6_12_r1;
    din_valid_6_13 <= out_new_pkt | hash_out_valid_filter_6_13;
    din_valid_6_13_r1 <= din_valid_6_13;
    din_valid_6_13_r2 <= din_valid_6_13_r1;

    din_6_13.data <= hash_out_valid_filter_6_13 ? hash_out_6_13 : 0;
    din_6_13.last <= out_new_pkt;
    din_6_13.bucket <= 6;


    din_6_13_r1 <= din_6_13;
    din_6_13_r2 <= din_6_13_r1;
    din_valid_6_14 <= out_new_pkt | hash_out_valid_filter_6_14;
    din_valid_6_14_r1 <= din_valid_6_14;
    din_valid_6_14_r2 <= din_valid_6_14_r1;

    din_6_14.data <= hash_out_valid_filter_6_14 ? hash_out_6_14 : 0;
    din_6_14.last <= out_new_pkt;
    din_6_14.bucket <= 6;


    din_6_14_r1 <= din_6_14;
    din_6_14_r2 <= din_6_14_r1;
    din_valid_6_15 <= out_new_pkt | hash_out_valid_filter_6_15;
    din_valid_6_15_r1 <= din_valid_6_15;
    din_valid_6_15_r2 <= din_valid_6_15_r1;

    din_6_15.data <= hash_out_valid_filter_6_15 ? hash_out_6_15 : 0;
    din_6_15.last <= out_new_pkt;
    din_6_15.bucket <= 6;


    din_6_15_r1 <= din_6_15;
    din_6_15_r2 <= din_6_15_r1;
    din_valid_6_16 <= out_new_pkt | hash_out_valid_filter_6_16;
    din_valid_6_16_r1 <= din_valid_6_16;
    din_valid_6_16_r2 <= din_valid_6_16_r1;

    din_6_16.data <= hash_out_valid_filter_6_16 ? hash_out_6_16 : 0;
    din_6_16.last <= out_new_pkt;
    din_6_16.bucket <= 6;


    din_6_16_r1 <= din_6_16;
    din_6_16_r2 <= din_6_16_r1;
    din_valid_6_17 <= out_new_pkt | hash_out_valid_filter_6_17;
    din_valid_6_17_r1 <= din_valid_6_17;
    din_valid_6_17_r2 <= din_valid_6_17_r1;

    din_6_17.data <= hash_out_valid_filter_6_17 ? hash_out_6_17 : 0;
    din_6_17.last <= out_new_pkt;
    din_6_17.bucket <= 6;


    din_6_17_r1 <= din_6_17;
    din_6_17_r2 <= din_6_17_r1;
    din_valid_6_18 <= out_new_pkt | hash_out_valid_filter_6_18;
    din_valid_6_18_r1 <= din_valid_6_18;
    din_valid_6_18_r2 <= din_valid_6_18_r1;

    din_6_18.data <= hash_out_valid_filter_6_18 ? hash_out_6_18 : 0;
    din_6_18.last <= out_new_pkt;
    din_6_18.bucket <= 6;


    din_6_18_r1 <= din_6_18;
    din_6_18_r2 <= din_6_18_r1;
    din_valid_6_19 <= out_new_pkt | hash_out_valid_filter_6_19;
    din_valid_6_19_r1 <= din_valid_6_19;
    din_valid_6_19_r2 <= din_valid_6_19_r1;

    din_6_19.data <= hash_out_valid_filter_6_19 ? hash_out_6_19 : 0;
    din_6_19.last <= out_new_pkt;
    din_6_19.bucket <= 6;


    din_6_19_r1 <= din_6_19;
    din_6_19_r2 <= din_6_19_r1;
    din_valid_6_20 <= out_new_pkt | hash_out_valid_filter_6_20;
    din_valid_6_20_r1 <= din_valid_6_20;
    din_valid_6_20_r2 <= din_valid_6_20_r1;

    din_6_20.data <= hash_out_valid_filter_6_20 ? hash_out_6_20 : 0;
    din_6_20.last <= out_new_pkt;
    din_6_20.bucket <= 6;


    din_6_20_r1 <= din_6_20;
    din_6_20_r2 <= din_6_20_r1;
    din_valid_6_21 <= out_new_pkt | hash_out_valid_filter_6_21;
    din_valid_6_21_r1 <= din_valid_6_21;
    din_valid_6_21_r2 <= din_valid_6_21_r1;

    din_6_21.data <= hash_out_valid_filter_6_21 ? hash_out_6_21 : 0;
    din_6_21.last <= out_new_pkt;
    din_6_21.bucket <= 6;


    din_6_21_r1 <= din_6_21;
    din_6_21_r2 <= din_6_21_r1;
    din_valid_6_22 <= out_new_pkt | hash_out_valid_filter_6_22;
    din_valid_6_22_r1 <= din_valid_6_22;
    din_valid_6_22_r2 <= din_valid_6_22_r1;

    din_6_22.data <= hash_out_valid_filter_6_22 ? hash_out_6_22 : 0;
    din_6_22.last <= out_new_pkt;
    din_6_22.bucket <= 6;


    din_6_22_r1 <= din_6_22;
    din_6_22_r2 <= din_6_22_r1;
    din_valid_6_23 <= out_new_pkt | hash_out_valid_filter_6_23;
    din_valid_6_23_r1 <= din_valid_6_23;
    din_valid_6_23_r2 <= din_valid_6_23_r1;

    din_6_23.data <= hash_out_valid_filter_6_23 ? hash_out_6_23 : 0;
    din_6_23.last <= out_new_pkt;
    din_6_23.bucket <= 6;


    din_6_23_r1 <= din_6_23;
    din_6_23_r2 <= din_6_23_r1;
    din_valid_6_24 <= out_new_pkt | hash_out_valid_filter_6_24;
    din_valid_6_24_r1 <= din_valid_6_24;
    din_valid_6_24_r2 <= din_valid_6_24_r1;

    din_6_24.data <= hash_out_valid_filter_6_24 ? hash_out_6_24 : 0;
    din_6_24.last <= out_new_pkt;
    din_6_24.bucket <= 6;


    din_6_24_r1 <= din_6_24;
    din_6_24_r2 <= din_6_24_r1;
    din_valid_6_25 <= out_new_pkt | hash_out_valid_filter_6_25;
    din_valid_6_25_r1 <= din_valid_6_25;
    din_valid_6_25_r2 <= din_valid_6_25_r1;

    din_6_25.data <= hash_out_valid_filter_6_25 ? hash_out_6_25 : 0;
    din_6_25.last <= out_new_pkt;
    din_6_25.bucket <= 6;


    din_6_25_r1 <= din_6_25;
    din_6_25_r2 <= din_6_25_r1;
    din_valid_6_26 <= out_new_pkt | hash_out_valid_filter_6_26;
    din_valid_6_26_r1 <= din_valid_6_26;
    din_valid_6_26_r2 <= din_valid_6_26_r1;

    din_6_26.data <= hash_out_valid_filter_6_26 ? hash_out_6_26 : 0;
    din_6_26.last <= out_new_pkt;
    din_6_26.bucket <= 6;


    din_6_26_r1 <= din_6_26;
    din_6_26_r2 <= din_6_26_r1;
    din_valid_6_27 <= out_new_pkt | hash_out_valid_filter_6_27;
    din_valid_6_27_r1 <= din_valid_6_27;
    din_valid_6_27_r2 <= din_valid_6_27_r1;

    din_6_27.data <= hash_out_valid_filter_6_27 ? hash_out_6_27 : 0;
    din_6_27.last <= out_new_pkt;
    din_6_27.bucket <= 6;


    din_6_27_r1 <= din_6_27;
    din_6_27_r2 <= din_6_27_r1;
    din_valid_6_28 <= out_new_pkt | hash_out_valid_filter_6_28;
    din_valid_6_28_r1 <= din_valid_6_28;
    din_valid_6_28_r2 <= din_valid_6_28_r1;

    din_6_28.data <= hash_out_valid_filter_6_28 ? hash_out_6_28 : 0;
    din_6_28.last <= out_new_pkt;
    din_6_28.bucket <= 6;


    din_6_28_r1 <= din_6_28;
    din_6_28_r2 <= din_6_28_r1;
    din_valid_6_29 <= out_new_pkt | hash_out_valid_filter_6_29;
    din_valid_6_29_r1 <= din_valid_6_29;
    din_valid_6_29_r2 <= din_valid_6_29_r1;

    din_6_29.data <= hash_out_valid_filter_6_29 ? hash_out_6_29 : 0;
    din_6_29.last <= out_new_pkt;
    din_6_29.bucket <= 6;


    din_6_29_r1 <= din_6_29;
    din_6_29_r2 <= din_6_29_r1;
    din_valid_6_30 <= out_new_pkt | hash_out_valid_filter_6_30;
    din_valid_6_30_r1 <= din_valid_6_30;
    din_valid_6_30_r2 <= din_valid_6_30_r1;

    din_6_30.data <= hash_out_valid_filter_6_30 ? hash_out_6_30 : 0;
    din_6_30.last <= out_new_pkt;
    din_6_30.bucket <= 6;


    din_6_30_r1 <= din_6_30;
    din_6_30_r2 <= din_6_30_r1;
    din_valid_6_31 <= out_new_pkt | hash_out_valid_filter_6_31;
    din_valid_6_31_r1 <= din_valid_6_31;
    din_valid_6_31_r2 <= din_valid_6_31_r1;

    din_6_31.data <= hash_out_valid_filter_6_31 ? hash_out_6_31 : 0;
    din_6_31.last <= out_new_pkt;
    din_6_31.bucket <= 6;


    din_6_31_r1 <= din_6_31;
    din_6_31_r2 <= din_6_31_r1;
    din_valid_7_0 <= out_new_pkt | hash_out_valid_filter_7_0;
    din_valid_7_0_r1 <= din_valid_7_0;
    din_valid_7_0_r2 <= din_valid_7_0_r1;

    din_7_0.data <= hash_out_valid_filter_7_0 ? hash_out_7_0 : 0;
    din_7_0.last <= out_new_pkt;
    din_7_0.bucket <= 7;


    din_7_0_r1 <= din_7_0;
    din_7_0_r2 <= din_7_0_r1;
    din_valid_7_1 <= out_new_pkt | hash_out_valid_filter_7_1;
    din_valid_7_1_r1 <= din_valid_7_1;
    din_valid_7_1_r2 <= din_valid_7_1_r1;

    din_7_1.data <= hash_out_valid_filter_7_1 ? hash_out_7_1 : 0;
    din_7_1.last <= out_new_pkt;
    din_7_1.bucket <= 7;


    din_7_1_r1 <= din_7_1;
    din_7_1_r2 <= din_7_1_r1;
    din_valid_7_2 <= out_new_pkt | hash_out_valid_filter_7_2;
    din_valid_7_2_r1 <= din_valid_7_2;
    din_valid_7_2_r2 <= din_valid_7_2_r1;

    din_7_2.data <= hash_out_valid_filter_7_2 ? hash_out_7_2 : 0;
    din_7_2.last <= out_new_pkt;
    din_7_2.bucket <= 7;


    din_7_2_r1 <= din_7_2;
    din_7_2_r2 <= din_7_2_r1;
    din_valid_7_3 <= out_new_pkt | hash_out_valid_filter_7_3;
    din_valid_7_3_r1 <= din_valid_7_3;
    din_valid_7_3_r2 <= din_valid_7_3_r1;

    din_7_3.data <= hash_out_valid_filter_7_3 ? hash_out_7_3 : 0;
    din_7_3.last <= out_new_pkt;
    din_7_3.bucket <= 7;


    din_7_3_r1 <= din_7_3;
    din_7_3_r2 <= din_7_3_r1;
    din_valid_7_4 <= out_new_pkt | hash_out_valid_filter_7_4;
    din_valid_7_4_r1 <= din_valid_7_4;
    din_valid_7_4_r2 <= din_valid_7_4_r1;

    din_7_4.data <= hash_out_valid_filter_7_4 ? hash_out_7_4 : 0;
    din_7_4.last <= out_new_pkt;
    din_7_4.bucket <= 7;


    din_7_4_r1 <= din_7_4;
    din_7_4_r2 <= din_7_4_r1;
    din_valid_7_5 <= out_new_pkt | hash_out_valid_filter_7_5;
    din_valid_7_5_r1 <= din_valid_7_5;
    din_valid_7_5_r2 <= din_valid_7_5_r1;

    din_7_5.data <= hash_out_valid_filter_7_5 ? hash_out_7_5 : 0;
    din_7_5.last <= out_new_pkt;
    din_7_5.bucket <= 7;


    din_7_5_r1 <= din_7_5;
    din_7_5_r2 <= din_7_5_r1;
    din_valid_7_6 <= out_new_pkt | hash_out_valid_filter_7_6;
    din_valid_7_6_r1 <= din_valid_7_6;
    din_valid_7_6_r2 <= din_valid_7_6_r1;

    din_7_6.data <= hash_out_valid_filter_7_6 ? hash_out_7_6 : 0;
    din_7_6.last <= out_new_pkt;
    din_7_6.bucket <= 7;


    din_7_6_r1 <= din_7_6;
    din_7_6_r2 <= din_7_6_r1;
    din_valid_7_7 <= out_new_pkt | hash_out_valid_filter_7_7;
    din_valid_7_7_r1 <= din_valid_7_7;
    din_valid_7_7_r2 <= din_valid_7_7_r1;

    din_7_7.data <= hash_out_valid_filter_7_7 ? hash_out_7_7 : 0;
    din_7_7.last <= out_new_pkt;
    din_7_7.bucket <= 7;


    din_7_7_r1 <= din_7_7;
    din_7_7_r2 <= din_7_7_r1;
    din_valid_7_8 <= out_new_pkt | hash_out_valid_filter_7_8;
    din_valid_7_8_r1 <= din_valid_7_8;
    din_valid_7_8_r2 <= din_valid_7_8_r1;

    din_7_8.data <= hash_out_valid_filter_7_8 ? hash_out_7_8 : 0;
    din_7_8.last <= out_new_pkt;
    din_7_8.bucket <= 7;


    din_7_8_r1 <= din_7_8;
    din_7_8_r2 <= din_7_8_r1;
    din_valid_7_9 <= out_new_pkt | hash_out_valid_filter_7_9;
    din_valid_7_9_r1 <= din_valid_7_9;
    din_valid_7_9_r2 <= din_valid_7_9_r1;

    din_7_9.data <= hash_out_valid_filter_7_9 ? hash_out_7_9 : 0;
    din_7_9.last <= out_new_pkt;
    din_7_9.bucket <= 7;


    din_7_9_r1 <= din_7_9;
    din_7_9_r2 <= din_7_9_r1;
    din_valid_7_10 <= out_new_pkt | hash_out_valid_filter_7_10;
    din_valid_7_10_r1 <= din_valid_7_10;
    din_valid_7_10_r2 <= din_valid_7_10_r1;

    din_7_10.data <= hash_out_valid_filter_7_10 ? hash_out_7_10 : 0;
    din_7_10.last <= out_new_pkt;
    din_7_10.bucket <= 7;


    din_7_10_r1 <= din_7_10;
    din_7_10_r2 <= din_7_10_r1;
    din_valid_7_11 <= out_new_pkt | hash_out_valid_filter_7_11;
    din_valid_7_11_r1 <= din_valid_7_11;
    din_valid_7_11_r2 <= din_valid_7_11_r1;

    din_7_11.data <= hash_out_valid_filter_7_11 ? hash_out_7_11 : 0;
    din_7_11.last <= out_new_pkt;
    din_7_11.bucket <= 7;


    din_7_11_r1 <= din_7_11;
    din_7_11_r2 <= din_7_11_r1;
    din_valid_7_12 <= out_new_pkt | hash_out_valid_filter_7_12;
    din_valid_7_12_r1 <= din_valid_7_12;
    din_valid_7_12_r2 <= din_valid_7_12_r1;

    din_7_12.data <= hash_out_valid_filter_7_12 ? hash_out_7_12 : 0;
    din_7_12.last <= out_new_pkt;
    din_7_12.bucket <= 7;


    din_7_12_r1 <= din_7_12;
    din_7_12_r2 <= din_7_12_r1;
    din_valid_7_13 <= out_new_pkt | hash_out_valid_filter_7_13;
    din_valid_7_13_r1 <= din_valid_7_13;
    din_valid_7_13_r2 <= din_valid_7_13_r1;

    din_7_13.data <= hash_out_valid_filter_7_13 ? hash_out_7_13 : 0;
    din_7_13.last <= out_new_pkt;
    din_7_13.bucket <= 7;


    din_7_13_r1 <= din_7_13;
    din_7_13_r2 <= din_7_13_r1;
    din_valid_7_14 <= out_new_pkt | hash_out_valid_filter_7_14;
    din_valid_7_14_r1 <= din_valid_7_14;
    din_valid_7_14_r2 <= din_valid_7_14_r1;

    din_7_14.data <= hash_out_valid_filter_7_14 ? hash_out_7_14 : 0;
    din_7_14.last <= out_new_pkt;
    din_7_14.bucket <= 7;


    din_7_14_r1 <= din_7_14;
    din_7_14_r2 <= din_7_14_r1;
    din_valid_7_15 <= out_new_pkt | hash_out_valid_filter_7_15;
    din_valid_7_15_r1 <= din_valid_7_15;
    din_valid_7_15_r2 <= din_valid_7_15_r1;

    din_7_15.data <= hash_out_valid_filter_7_15 ? hash_out_7_15 : 0;
    din_7_15.last <= out_new_pkt;
    din_7_15.bucket <= 7;


    din_7_15_r1 <= din_7_15;
    din_7_15_r2 <= din_7_15_r1;
    din_valid_7_16 <= out_new_pkt | hash_out_valid_filter_7_16;
    din_valid_7_16_r1 <= din_valid_7_16;
    din_valid_7_16_r2 <= din_valid_7_16_r1;

    din_7_16.data <= hash_out_valid_filter_7_16 ? hash_out_7_16 : 0;
    din_7_16.last <= out_new_pkt;
    din_7_16.bucket <= 7;


    din_7_16_r1 <= din_7_16;
    din_7_16_r2 <= din_7_16_r1;
    din_valid_7_17 <= out_new_pkt | hash_out_valid_filter_7_17;
    din_valid_7_17_r1 <= din_valid_7_17;
    din_valid_7_17_r2 <= din_valid_7_17_r1;

    din_7_17.data <= hash_out_valid_filter_7_17 ? hash_out_7_17 : 0;
    din_7_17.last <= out_new_pkt;
    din_7_17.bucket <= 7;


    din_7_17_r1 <= din_7_17;
    din_7_17_r2 <= din_7_17_r1;
    din_valid_7_18 <= out_new_pkt | hash_out_valid_filter_7_18;
    din_valid_7_18_r1 <= din_valid_7_18;
    din_valid_7_18_r2 <= din_valid_7_18_r1;

    din_7_18.data <= hash_out_valid_filter_7_18 ? hash_out_7_18 : 0;
    din_7_18.last <= out_new_pkt;
    din_7_18.bucket <= 7;


    din_7_18_r1 <= din_7_18;
    din_7_18_r2 <= din_7_18_r1;
    din_valid_7_19 <= out_new_pkt | hash_out_valid_filter_7_19;
    din_valid_7_19_r1 <= din_valid_7_19;
    din_valid_7_19_r2 <= din_valid_7_19_r1;

    din_7_19.data <= hash_out_valid_filter_7_19 ? hash_out_7_19 : 0;
    din_7_19.last <= out_new_pkt;
    din_7_19.bucket <= 7;


    din_7_19_r1 <= din_7_19;
    din_7_19_r2 <= din_7_19_r1;
    din_valid_7_20 <= out_new_pkt | hash_out_valid_filter_7_20;
    din_valid_7_20_r1 <= din_valid_7_20;
    din_valid_7_20_r2 <= din_valid_7_20_r1;

    din_7_20.data <= hash_out_valid_filter_7_20 ? hash_out_7_20 : 0;
    din_7_20.last <= out_new_pkt;
    din_7_20.bucket <= 7;


    din_7_20_r1 <= din_7_20;
    din_7_20_r2 <= din_7_20_r1;
    din_valid_7_21 <= out_new_pkt | hash_out_valid_filter_7_21;
    din_valid_7_21_r1 <= din_valid_7_21;
    din_valid_7_21_r2 <= din_valid_7_21_r1;

    din_7_21.data <= hash_out_valid_filter_7_21 ? hash_out_7_21 : 0;
    din_7_21.last <= out_new_pkt;
    din_7_21.bucket <= 7;


    din_7_21_r1 <= din_7_21;
    din_7_21_r2 <= din_7_21_r1;
    din_valid_7_22 <= out_new_pkt | hash_out_valid_filter_7_22;
    din_valid_7_22_r1 <= din_valid_7_22;
    din_valid_7_22_r2 <= din_valid_7_22_r1;

    din_7_22.data <= hash_out_valid_filter_7_22 ? hash_out_7_22 : 0;
    din_7_22.last <= out_new_pkt;
    din_7_22.bucket <= 7;


    din_7_22_r1 <= din_7_22;
    din_7_22_r2 <= din_7_22_r1;
    din_valid_7_23 <= out_new_pkt | hash_out_valid_filter_7_23;
    din_valid_7_23_r1 <= din_valid_7_23;
    din_valid_7_23_r2 <= din_valid_7_23_r1;

    din_7_23.data <= hash_out_valid_filter_7_23 ? hash_out_7_23 : 0;
    din_7_23.last <= out_new_pkt;
    din_7_23.bucket <= 7;


    din_7_23_r1 <= din_7_23;
    din_7_23_r2 <= din_7_23_r1;
    din_valid_7_24 <= out_new_pkt | hash_out_valid_filter_7_24;
    din_valid_7_24_r1 <= din_valid_7_24;
    din_valid_7_24_r2 <= din_valid_7_24_r1;

    din_7_24.data <= hash_out_valid_filter_7_24 ? hash_out_7_24 : 0;
    din_7_24.last <= out_new_pkt;
    din_7_24.bucket <= 7;


    din_7_24_r1 <= din_7_24;
    din_7_24_r2 <= din_7_24_r1;
    din_valid_7_25 <= out_new_pkt | hash_out_valid_filter_7_25;
    din_valid_7_25_r1 <= din_valid_7_25;
    din_valid_7_25_r2 <= din_valid_7_25_r1;

    din_7_25.data <= hash_out_valid_filter_7_25 ? hash_out_7_25 : 0;
    din_7_25.last <= out_new_pkt;
    din_7_25.bucket <= 7;


    din_7_25_r1 <= din_7_25;
    din_7_25_r2 <= din_7_25_r1;
    din_valid_7_26 <= out_new_pkt | hash_out_valid_filter_7_26;
    din_valid_7_26_r1 <= din_valid_7_26;
    din_valid_7_26_r2 <= din_valid_7_26_r1;

    din_7_26.data <= hash_out_valid_filter_7_26 ? hash_out_7_26 : 0;
    din_7_26.last <= out_new_pkt;
    din_7_26.bucket <= 7;


    din_7_26_r1 <= din_7_26;
    din_7_26_r2 <= din_7_26_r1;
    din_valid_7_27 <= out_new_pkt | hash_out_valid_filter_7_27;
    din_valid_7_27_r1 <= din_valid_7_27;
    din_valid_7_27_r2 <= din_valid_7_27_r1;

    din_7_27.data <= hash_out_valid_filter_7_27 ? hash_out_7_27 : 0;
    din_7_27.last <= out_new_pkt;
    din_7_27.bucket <= 7;


    din_7_27_r1 <= din_7_27;
    din_7_27_r2 <= din_7_27_r1;
    din_valid_7_28 <= out_new_pkt | hash_out_valid_filter_7_28;
    din_valid_7_28_r1 <= din_valid_7_28;
    din_valid_7_28_r2 <= din_valid_7_28_r1;

    din_7_28.data <= hash_out_valid_filter_7_28 ? hash_out_7_28 : 0;
    din_7_28.last <= out_new_pkt;
    din_7_28.bucket <= 7;


    din_7_28_r1 <= din_7_28;
    din_7_28_r2 <= din_7_28_r1;
    din_valid_7_29 <= out_new_pkt | hash_out_valid_filter_7_29;
    din_valid_7_29_r1 <= din_valid_7_29;
    din_valid_7_29_r2 <= din_valid_7_29_r1;

    din_7_29.data <= hash_out_valid_filter_7_29 ? hash_out_7_29 : 0;
    din_7_29.last <= out_new_pkt;
    din_7_29.bucket <= 7;


    din_7_29_r1 <= din_7_29;
    din_7_29_r2 <= din_7_29_r1;
    din_valid_7_30 <= out_new_pkt | hash_out_valid_filter_7_30;
    din_valid_7_30_r1 <= din_valid_7_30;
    din_valid_7_30_r2 <= din_valid_7_30_r1;

    din_7_30.data <= hash_out_valid_filter_7_30 ? hash_out_7_30 : 0;
    din_7_30.last <= out_new_pkt;
    din_7_30.bucket <= 7;


    din_7_30_r1 <= din_7_30;
    din_7_30_r2 <= din_7_30_r1;
    din_valid_7_31 <= out_new_pkt | hash_out_valid_filter_7_31;
    din_valid_7_31_r1 <= din_valid_7_31;
    din_valid_7_31_r2 <= din_valid_7_31_r1;

    din_7_31.data <= hash_out_valid_filter_7_31 ? hash_out_7_31 : 0;
    din_7_31.last <= out_new_pkt;
    din_7_31.bucket <= 7;


    din_7_31_r1 <= din_7_31;
    din_7_31_r2 <= din_7_31_r1;
end

//Instantiation
simple_fifo #(
    .DATA_WIDTH(META_WIDTH),
    .ADDR_WIDTH(9)
) meta_fifo (
	.clk               (clk),                      
	.rst               (rst),            
	.din               (in_meta_data),          
	.din_valid         (in_meta_valid),         
	.din_ready         (in_meta_ready),         
	.dout              (internal_meta_data),                        
	.dout_valid        (internal_meta_valid),                       
	.dout_ready        (internal_meta_ready)                       
);


frontend front(
    .clk(clk),
    .rst(rst),
    .hash_out_0_0(hash_out_0_0),
    .hash_out_valid_filter_0_0(hash_out_valid_filter_0_0),
    .hash_out_0_1(hash_out_0_1),
    .hash_out_valid_filter_0_1(hash_out_valid_filter_0_1),
    .hash_out_0_2(hash_out_0_2),
    .hash_out_valid_filter_0_2(hash_out_valid_filter_0_2),
    .hash_out_0_3(hash_out_0_3),
    .hash_out_valid_filter_0_3(hash_out_valid_filter_0_3),
    .hash_out_0_4(hash_out_0_4),
    .hash_out_valid_filter_0_4(hash_out_valid_filter_0_4),
    .hash_out_0_5(hash_out_0_5),
    .hash_out_valid_filter_0_5(hash_out_valid_filter_0_5),
    .hash_out_0_6(hash_out_0_6),
    .hash_out_valid_filter_0_6(hash_out_valid_filter_0_6),
    .hash_out_0_7(hash_out_0_7),
    .hash_out_valid_filter_0_7(hash_out_valid_filter_0_7),
    .hash_out_0_8(hash_out_0_8),
    .hash_out_valid_filter_0_8(hash_out_valid_filter_0_8),
    .hash_out_0_9(hash_out_0_9),
    .hash_out_valid_filter_0_9(hash_out_valid_filter_0_9),
    .hash_out_0_10(hash_out_0_10),
    .hash_out_valid_filter_0_10(hash_out_valid_filter_0_10),
    .hash_out_0_11(hash_out_0_11),
    .hash_out_valid_filter_0_11(hash_out_valid_filter_0_11),
    .hash_out_0_12(hash_out_0_12),
    .hash_out_valid_filter_0_12(hash_out_valid_filter_0_12),
    .hash_out_0_13(hash_out_0_13),
    .hash_out_valid_filter_0_13(hash_out_valid_filter_0_13),
    .hash_out_0_14(hash_out_0_14),
    .hash_out_valid_filter_0_14(hash_out_valid_filter_0_14),
    .hash_out_0_15(hash_out_0_15),
    .hash_out_valid_filter_0_15(hash_out_valid_filter_0_15),
    .hash_out_0_16(hash_out_0_16),
    .hash_out_valid_filter_0_16(hash_out_valid_filter_0_16),
    .hash_out_0_17(hash_out_0_17),
    .hash_out_valid_filter_0_17(hash_out_valid_filter_0_17),
    .hash_out_0_18(hash_out_0_18),
    .hash_out_valid_filter_0_18(hash_out_valid_filter_0_18),
    .hash_out_0_19(hash_out_0_19),
    .hash_out_valid_filter_0_19(hash_out_valid_filter_0_19),
    .hash_out_0_20(hash_out_0_20),
    .hash_out_valid_filter_0_20(hash_out_valid_filter_0_20),
    .hash_out_0_21(hash_out_0_21),
    .hash_out_valid_filter_0_21(hash_out_valid_filter_0_21),
    .hash_out_0_22(hash_out_0_22),
    .hash_out_valid_filter_0_22(hash_out_valid_filter_0_22),
    .hash_out_0_23(hash_out_0_23),
    .hash_out_valid_filter_0_23(hash_out_valid_filter_0_23),
    .hash_out_0_24(hash_out_0_24),
    .hash_out_valid_filter_0_24(hash_out_valid_filter_0_24),
    .hash_out_0_25(hash_out_0_25),
    .hash_out_valid_filter_0_25(hash_out_valid_filter_0_25),
    .hash_out_0_26(hash_out_0_26),
    .hash_out_valid_filter_0_26(hash_out_valid_filter_0_26),
    .hash_out_0_27(hash_out_0_27),
    .hash_out_valid_filter_0_27(hash_out_valid_filter_0_27),
    .hash_out_0_28(hash_out_0_28),
    .hash_out_valid_filter_0_28(hash_out_valid_filter_0_28),
    .hash_out_0_29(hash_out_0_29),
    .hash_out_valid_filter_0_29(hash_out_valid_filter_0_29),
    .hash_out_0_30(hash_out_0_30),
    .hash_out_valid_filter_0_30(hash_out_valid_filter_0_30),
    .hash_out_0_31(hash_out_0_31),
    .hash_out_valid_filter_0_31(hash_out_valid_filter_0_31),
    .hash_out_1_0(hash_out_1_0),
    .hash_out_valid_filter_1_0(hash_out_valid_filter_1_0),
    .hash_out_1_1(hash_out_1_1),
    .hash_out_valid_filter_1_1(hash_out_valid_filter_1_1),
    .hash_out_1_2(hash_out_1_2),
    .hash_out_valid_filter_1_2(hash_out_valid_filter_1_2),
    .hash_out_1_3(hash_out_1_3),
    .hash_out_valid_filter_1_3(hash_out_valid_filter_1_3),
    .hash_out_1_4(hash_out_1_4),
    .hash_out_valid_filter_1_4(hash_out_valid_filter_1_4),
    .hash_out_1_5(hash_out_1_5),
    .hash_out_valid_filter_1_5(hash_out_valid_filter_1_5),
    .hash_out_1_6(hash_out_1_6),
    .hash_out_valid_filter_1_6(hash_out_valid_filter_1_6),
    .hash_out_1_7(hash_out_1_7),
    .hash_out_valid_filter_1_7(hash_out_valid_filter_1_7),
    .hash_out_1_8(hash_out_1_8),
    .hash_out_valid_filter_1_8(hash_out_valid_filter_1_8),
    .hash_out_1_9(hash_out_1_9),
    .hash_out_valid_filter_1_9(hash_out_valid_filter_1_9),
    .hash_out_1_10(hash_out_1_10),
    .hash_out_valid_filter_1_10(hash_out_valid_filter_1_10),
    .hash_out_1_11(hash_out_1_11),
    .hash_out_valid_filter_1_11(hash_out_valid_filter_1_11),
    .hash_out_1_12(hash_out_1_12),
    .hash_out_valid_filter_1_12(hash_out_valid_filter_1_12),
    .hash_out_1_13(hash_out_1_13),
    .hash_out_valid_filter_1_13(hash_out_valid_filter_1_13),
    .hash_out_1_14(hash_out_1_14),
    .hash_out_valid_filter_1_14(hash_out_valid_filter_1_14),
    .hash_out_1_15(hash_out_1_15),
    .hash_out_valid_filter_1_15(hash_out_valid_filter_1_15),
    .hash_out_1_16(hash_out_1_16),
    .hash_out_valid_filter_1_16(hash_out_valid_filter_1_16),
    .hash_out_1_17(hash_out_1_17),
    .hash_out_valid_filter_1_17(hash_out_valid_filter_1_17),
    .hash_out_1_18(hash_out_1_18),
    .hash_out_valid_filter_1_18(hash_out_valid_filter_1_18),
    .hash_out_1_19(hash_out_1_19),
    .hash_out_valid_filter_1_19(hash_out_valid_filter_1_19),
    .hash_out_1_20(hash_out_1_20),
    .hash_out_valid_filter_1_20(hash_out_valid_filter_1_20),
    .hash_out_1_21(hash_out_1_21),
    .hash_out_valid_filter_1_21(hash_out_valid_filter_1_21),
    .hash_out_1_22(hash_out_1_22),
    .hash_out_valid_filter_1_22(hash_out_valid_filter_1_22),
    .hash_out_1_23(hash_out_1_23),
    .hash_out_valid_filter_1_23(hash_out_valid_filter_1_23),
    .hash_out_1_24(hash_out_1_24),
    .hash_out_valid_filter_1_24(hash_out_valid_filter_1_24),
    .hash_out_1_25(hash_out_1_25),
    .hash_out_valid_filter_1_25(hash_out_valid_filter_1_25),
    .hash_out_1_26(hash_out_1_26),
    .hash_out_valid_filter_1_26(hash_out_valid_filter_1_26),
    .hash_out_1_27(hash_out_1_27),
    .hash_out_valid_filter_1_27(hash_out_valid_filter_1_27),
    .hash_out_1_28(hash_out_1_28),
    .hash_out_valid_filter_1_28(hash_out_valid_filter_1_28),
    .hash_out_1_29(hash_out_1_29),
    .hash_out_valid_filter_1_29(hash_out_valid_filter_1_29),
    .hash_out_1_30(hash_out_1_30),
    .hash_out_valid_filter_1_30(hash_out_valid_filter_1_30),
    .hash_out_1_31(hash_out_1_31),
    .hash_out_valid_filter_1_31(hash_out_valid_filter_1_31),
    .hash_out_2_0(hash_out_2_0),
    .hash_out_valid_filter_2_0(hash_out_valid_filter_2_0),
    .hash_out_2_1(hash_out_2_1),
    .hash_out_valid_filter_2_1(hash_out_valid_filter_2_1),
    .hash_out_2_2(hash_out_2_2),
    .hash_out_valid_filter_2_2(hash_out_valid_filter_2_2),
    .hash_out_2_3(hash_out_2_3),
    .hash_out_valid_filter_2_3(hash_out_valid_filter_2_3),
    .hash_out_2_4(hash_out_2_4),
    .hash_out_valid_filter_2_4(hash_out_valid_filter_2_4),
    .hash_out_2_5(hash_out_2_5),
    .hash_out_valid_filter_2_5(hash_out_valid_filter_2_5),
    .hash_out_2_6(hash_out_2_6),
    .hash_out_valid_filter_2_6(hash_out_valid_filter_2_6),
    .hash_out_2_7(hash_out_2_7),
    .hash_out_valid_filter_2_7(hash_out_valid_filter_2_7),
    .hash_out_2_8(hash_out_2_8),
    .hash_out_valid_filter_2_8(hash_out_valid_filter_2_8),
    .hash_out_2_9(hash_out_2_9),
    .hash_out_valid_filter_2_9(hash_out_valid_filter_2_9),
    .hash_out_2_10(hash_out_2_10),
    .hash_out_valid_filter_2_10(hash_out_valid_filter_2_10),
    .hash_out_2_11(hash_out_2_11),
    .hash_out_valid_filter_2_11(hash_out_valid_filter_2_11),
    .hash_out_2_12(hash_out_2_12),
    .hash_out_valid_filter_2_12(hash_out_valid_filter_2_12),
    .hash_out_2_13(hash_out_2_13),
    .hash_out_valid_filter_2_13(hash_out_valid_filter_2_13),
    .hash_out_2_14(hash_out_2_14),
    .hash_out_valid_filter_2_14(hash_out_valid_filter_2_14),
    .hash_out_2_15(hash_out_2_15),
    .hash_out_valid_filter_2_15(hash_out_valid_filter_2_15),
    .hash_out_2_16(hash_out_2_16),
    .hash_out_valid_filter_2_16(hash_out_valid_filter_2_16),
    .hash_out_2_17(hash_out_2_17),
    .hash_out_valid_filter_2_17(hash_out_valid_filter_2_17),
    .hash_out_2_18(hash_out_2_18),
    .hash_out_valid_filter_2_18(hash_out_valid_filter_2_18),
    .hash_out_2_19(hash_out_2_19),
    .hash_out_valid_filter_2_19(hash_out_valid_filter_2_19),
    .hash_out_2_20(hash_out_2_20),
    .hash_out_valid_filter_2_20(hash_out_valid_filter_2_20),
    .hash_out_2_21(hash_out_2_21),
    .hash_out_valid_filter_2_21(hash_out_valid_filter_2_21),
    .hash_out_2_22(hash_out_2_22),
    .hash_out_valid_filter_2_22(hash_out_valid_filter_2_22),
    .hash_out_2_23(hash_out_2_23),
    .hash_out_valid_filter_2_23(hash_out_valid_filter_2_23),
    .hash_out_2_24(hash_out_2_24),
    .hash_out_valid_filter_2_24(hash_out_valid_filter_2_24),
    .hash_out_2_25(hash_out_2_25),
    .hash_out_valid_filter_2_25(hash_out_valid_filter_2_25),
    .hash_out_2_26(hash_out_2_26),
    .hash_out_valid_filter_2_26(hash_out_valid_filter_2_26),
    .hash_out_2_27(hash_out_2_27),
    .hash_out_valid_filter_2_27(hash_out_valid_filter_2_27),
    .hash_out_2_28(hash_out_2_28),
    .hash_out_valid_filter_2_28(hash_out_valid_filter_2_28),
    .hash_out_2_29(hash_out_2_29),
    .hash_out_valid_filter_2_29(hash_out_valid_filter_2_29),
    .hash_out_2_30(hash_out_2_30),
    .hash_out_valid_filter_2_30(hash_out_valid_filter_2_30),
    .hash_out_2_31(hash_out_2_31),
    .hash_out_valid_filter_2_31(hash_out_valid_filter_2_31),
    .hash_out_3_0(hash_out_3_0),
    .hash_out_valid_filter_3_0(hash_out_valid_filter_3_0),
    .hash_out_3_1(hash_out_3_1),
    .hash_out_valid_filter_3_1(hash_out_valid_filter_3_1),
    .hash_out_3_2(hash_out_3_2),
    .hash_out_valid_filter_3_2(hash_out_valid_filter_3_2),
    .hash_out_3_3(hash_out_3_3),
    .hash_out_valid_filter_3_3(hash_out_valid_filter_3_3),
    .hash_out_3_4(hash_out_3_4),
    .hash_out_valid_filter_3_4(hash_out_valid_filter_3_4),
    .hash_out_3_5(hash_out_3_5),
    .hash_out_valid_filter_3_5(hash_out_valid_filter_3_5),
    .hash_out_3_6(hash_out_3_6),
    .hash_out_valid_filter_3_6(hash_out_valid_filter_3_6),
    .hash_out_3_7(hash_out_3_7),
    .hash_out_valid_filter_3_7(hash_out_valid_filter_3_7),
    .hash_out_3_8(hash_out_3_8),
    .hash_out_valid_filter_3_8(hash_out_valid_filter_3_8),
    .hash_out_3_9(hash_out_3_9),
    .hash_out_valid_filter_3_9(hash_out_valid_filter_3_9),
    .hash_out_3_10(hash_out_3_10),
    .hash_out_valid_filter_3_10(hash_out_valid_filter_3_10),
    .hash_out_3_11(hash_out_3_11),
    .hash_out_valid_filter_3_11(hash_out_valid_filter_3_11),
    .hash_out_3_12(hash_out_3_12),
    .hash_out_valid_filter_3_12(hash_out_valid_filter_3_12),
    .hash_out_3_13(hash_out_3_13),
    .hash_out_valid_filter_3_13(hash_out_valid_filter_3_13),
    .hash_out_3_14(hash_out_3_14),
    .hash_out_valid_filter_3_14(hash_out_valid_filter_3_14),
    .hash_out_3_15(hash_out_3_15),
    .hash_out_valid_filter_3_15(hash_out_valid_filter_3_15),
    .hash_out_3_16(hash_out_3_16),
    .hash_out_valid_filter_3_16(hash_out_valid_filter_3_16),
    .hash_out_3_17(hash_out_3_17),
    .hash_out_valid_filter_3_17(hash_out_valid_filter_3_17),
    .hash_out_3_18(hash_out_3_18),
    .hash_out_valid_filter_3_18(hash_out_valid_filter_3_18),
    .hash_out_3_19(hash_out_3_19),
    .hash_out_valid_filter_3_19(hash_out_valid_filter_3_19),
    .hash_out_3_20(hash_out_3_20),
    .hash_out_valid_filter_3_20(hash_out_valid_filter_3_20),
    .hash_out_3_21(hash_out_3_21),
    .hash_out_valid_filter_3_21(hash_out_valid_filter_3_21),
    .hash_out_3_22(hash_out_3_22),
    .hash_out_valid_filter_3_22(hash_out_valid_filter_3_22),
    .hash_out_3_23(hash_out_3_23),
    .hash_out_valid_filter_3_23(hash_out_valid_filter_3_23),
    .hash_out_3_24(hash_out_3_24),
    .hash_out_valid_filter_3_24(hash_out_valid_filter_3_24),
    .hash_out_3_25(hash_out_3_25),
    .hash_out_valid_filter_3_25(hash_out_valid_filter_3_25),
    .hash_out_3_26(hash_out_3_26),
    .hash_out_valid_filter_3_26(hash_out_valid_filter_3_26),
    .hash_out_3_27(hash_out_3_27),
    .hash_out_valid_filter_3_27(hash_out_valid_filter_3_27),
    .hash_out_3_28(hash_out_3_28),
    .hash_out_valid_filter_3_28(hash_out_valid_filter_3_28),
    .hash_out_3_29(hash_out_3_29),
    .hash_out_valid_filter_3_29(hash_out_valid_filter_3_29),
    .hash_out_3_30(hash_out_3_30),
    .hash_out_valid_filter_3_30(hash_out_valid_filter_3_30),
    .hash_out_3_31(hash_out_3_31),
    .hash_out_valid_filter_3_31(hash_out_valid_filter_3_31),
    .hash_out_4_0(hash_out_4_0),
    .hash_out_valid_filter_4_0(hash_out_valid_filter_4_0),
    .hash_out_4_1(hash_out_4_1),
    .hash_out_valid_filter_4_1(hash_out_valid_filter_4_1),
    .hash_out_4_2(hash_out_4_2),
    .hash_out_valid_filter_4_2(hash_out_valid_filter_4_2),
    .hash_out_4_3(hash_out_4_3),
    .hash_out_valid_filter_4_3(hash_out_valid_filter_4_3),
    .hash_out_4_4(hash_out_4_4),
    .hash_out_valid_filter_4_4(hash_out_valid_filter_4_4),
    .hash_out_4_5(hash_out_4_5),
    .hash_out_valid_filter_4_5(hash_out_valid_filter_4_5),
    .hash_out_4_6(hash_out_4_6),
    .hash_out_valid_filter_4_6(hash_out_valid_filter_4_6),
    .hash_out_4_7(hash_out_4_7),
    .hash_out_valid_filter_4_7(hash_out_valid_filter_4_7),
    .hash_out_4_8(hash_out_4_8),
    .hash_out_valid_filter_4_8(hash_out_valid_filter_4_8),
    .hash_out_4_9(hash_out_4_9),
    .hash_out_valid_filter_4_9(hash_out_valid_filter_4_9),
    .hash_out_4_10(hash_out_4_10),
    .hash_out_valid_filter_4_10(hash_out_valid_filter_4_10),
    .hash_out_4_11(hash_out_4_11),
    .hash_out_valid_filter_4_11(hash_out_valid_filter_4_11),
    .hash_out_4_12(hash_out_4_12),
    .hash_out_valid_filter_4_12(hash_out_valid_filter_4_12),
    .hash_out_4_13(hash_out_4_13),
    .hash_out_valid_filter_4_13(hash_out_valid_filter_4_13),
    .hash_out_4_14(hash_out_4_14),
    .hash_out_valid_filter_4_14(hash_out_valid_filter_4_14),
    .hash_out_4_15(hash_out_4_15),
    .hash_out_valid_filter_4_15(hash_out_valid_filter_4_15),
    .hash_out_4_16(hash_out_4_16),
    .hash_out_valid_filter_4_16(hash_out_valid_filter_4_16),
    .hash_out_4_17(hash_out_4_17),
    .hash_out_valid_filter_4_17(hash_out_valid_filter_4_17),
    .hash_out_4_18(hash_out_4_18),
    .hash_out_valid_filter_4_18(hash_out_valid_filter_4_18),
    .hash_out_4_19(hash_out_4_19),
    .hash_out_valid_filter_4_19(hash_out_valid_filter_4_19),
    .hash_out_4_20(hash_out_4_20),
    .hash_out_valid_filter_4_20(hash_out_valid_filter_4_20),
    .hash_out_4_21(hash_out_4_21),
    .hash_out_valid_filter_4_21(hash_out_valid_filter_4_21),
    .hash_out_4_22(hash_out_4_22),
    .hash_out_valid_filter_4_22(hash_out_valid_filter_4_22),
    .hash_out_4_23(hash_out_4_23),
    .hash_out_valid_filter_4_23(hash_out_valid_filter_4_23),
    .hash_out_4_24(hash_out_4_24),
    .hash_out_valid_filter_4_24(hash_out_valid_filter_4_24),
    .hash_out_4_25(hash_out_4_25),
    .hash_out_valid_filter_4_25(hash_out_valid_filter_4_25),
    .hash_out_4_26(hash_out_4_26),
    .hash_out_valid_filter_4_26(hash_out_valid_filter_4_26),
    .hash_out_4_27(hash_out_4_27),
    .hash_out_valid_filter_4_27(hash_out_valid_filter_4_27),
    .hash_out_4_28(hash_out_4_28),
    .hash_out_valid_filter_4_28(hash_out_valid_filter_4_28),
    .hash_out_4_29(hash_out_4_29),
    .hash_out_valid_filter_4_29(hash_out_valid_filter_4_29),
    .hash_out_4_30(hash_out_4_30),
    .hash_out_valid_filter_4_30(hash_out_valid_filter_4_30),
    .hash_out_4_31(hash_out_4_31),
    .hash_out_valid_filter_4_31(hash_out_valid_filter_4_31),
    .hash_out_5_0(hash_out_5_0),
    .hash_out_valid_filter_5_0(hash_out_valid_filter_5_0),
    .hash_out_5_1(hash_out_5_1),
    .hash_out_valid_filter_5_1(hash_out_valid_filter_5_1),
    .hash_out_5_2(hash_out_5_2),
    .hash_out_valid_filter_5_2(hash_out_valid_filter_5_2),
    .hash_out_5_3(hash_out_5_3),
    .hash_out_valid_filter_5_3(hash_out_valid_filter_5_3),
    .hash_out_5_4(hash_out_5_4),
    .hash_out_valid_filter_5_4(hash_out_valid_filter_5_4),
    .hash_out_5_5(hash_out_5_5),
    .hash_out_valid_filter_5_5(hash_out_valid_filter_5_5),
    .hash_out_5_6(hash_out_5_6),
    .hash_out_valid_filter_5_6(hash_out_valid_filter_5_6),
    .hash_out_5_7(hash_out_5_7),
    .hash_out_valid_filter_5_7(hash_out_valid_filter_5_7),
    .hash_out_5_8(hash_out_5_8),
    .hash_out_valid_filter_5_8(hash_out_valid_filter_5_8),
    .hash_out_5_9(hash_out_5_9),
    .hash_out_valid_filter_5_9(hash_out_valid_filter_5_9),
    .hash_out_5_10(hash_out_5_10),
    .hash_out_valid_filter_5_10(hash_out_valid_filter_5_10),
    .hash_out_5_11(hash_out_5_11),
    .hash_out_valid_filter_5_11(hash_out_valid_filter_5_11),
    .hash_out_5_12(hash_out_5_12),
    .hash_out_valid_filter_5_12(hash_out_valid_filter_5_12),
    .hash_out_5_13(hash_out_5_13),
    .hash_out_valid_filter_5_13(hash_out_valid_filter_5_13),
    .hash_out_5_14(hash_out_5_14),
    .hash_out_valid_filter_5_14(hash_out_valid_filter_5_14),
    .hash_out_5_15(hash_out_5_15),
    .hash_out_valid_filter_5_15(hash_out_valid_filter_5_15),
    .hash_out_5_16(hash_out_5_16),
    .hash_out_valid_filter_5_16(hash_out_valid_filter_5_16),
    .hash_out_5_17(hash_out_5_17),
    .hash_out_valid_filter_5_17(hash_out_valid_filter_5_17),
    .hash_out_5_18(hash_out_5_18),
    .hash_out_valid_filter_5_18(hash_out_valid_filter_5_18),
    .hash_out_5_19(hash_out_5_19),
    .hash_out_valid_filter_5_19(hash_out_valid_filter_5_19),
    .hash_out_5_20(hash_out_5_20),
    .hash_out_valid_filter_5_20(hash_out_valid_filter_5_20),
    .hash_out_5_21(hash_out_5_21),
    .hash_out_valid_filter_5_21(hash_out_valid_filter_5_21),
    .hash_out_5_22(hash_out_5_22),
    .hash_out_valid_filter_5_22(hash_out_valid_filter_5_22),
    .hash_out_5_23(hash_out_5_23),
    .hash_out_valid_filter_5_23(hash_out_valid_filter_5_23),
    .hash_out_5_24(hash_out_5_24),
    .hash_out_valid_filter_5_24(hash_out_valid_filter_5_24),
    .hash_out_5_25(hash_out_5_25),
    .hash_out_valid_filter_5_25(hash_out_valid_filter_5_25),
    .hash_out_5_26(hash_out_5_26),
    .hash_out_valid_filter_5_26(hash_out_valid_filter_5_26),
    .hash_out_5_27(hash_out_5_27),
    .hash_out_valid_filter_5_27(hash_out_valid_filter_5_27),
    .hash_out_5_28(hash_out_5_28),
    .hash_out_valid_filter_5_28(hash_out_valid_filter_5_28),
    .hash_out_5_29(hash_out_5_29),
    .hash_out_valid_filter_5_29(hash_out_valid_filter_5_29),
    .hash_out_5_30(hash_out_5_30),
    .hash_out_valid_filter_5_30(hash_out_valid_filter_5_30),
    .hash_out_5_31(hash_out_5_31),
    .hash_out_valid_filter_5_31(hash_out_valid_filter_5_31),
    .hash_out_6_0(hash_out_6_0),
    .hash_out_valid_filter_6_0(hash_out_valid_filter_6_0),
    .hash_out_6_1(hash_out_6_1),
    .hash_out_valid_filter_6_1(hash_out_valid_filter_6_1),
    .hash_out_6_2(hash_out_6_2),
    .hash_out_valid_filter_6_2(hash_out_valid_filter_6_2),
    .hash_out_6_3(hash_out_6_3),
    .hash_out_valid_filter_6_3(hash_out_valid_filter_6_3),
    .hash_out_6_4(hash_out_6_4),
    .hash_out_valid_filter_6_4(hash_out_valid_filter_6_4),
    .hash_out_6_5(hash_out_6_5),
    .hash_out_valid_filter_6_5(hash_out_valid_filter_6_5),
    .hash_out_6_6(hash_out_6_6),
    .hash_out_valid_filter_6_6(hash_out_valid_filter_6_6),
    .hash_out_6_7(hash_out_6_7),
    .hash_out_valid_filter_6_7(hash_out_valid_filter_6_7),
    .hash_out_6_8(hash_out_6_8),
    .hash_out_valid_filter_6_8(hash_out_valid_filter_6_8),
    .hash_out_6_9(hash_out_6_9),
    .hash_out_valid_filter_6_9(hash_out_valid_filter_6_9),
    .hash_out_6_10(hash_out_6_10),
    .hash_out_valid_filter_6_10(hash_out_valid_filter_6_10),
    .hash_out_6_11(hash_out_6_11),
    .hash_out_valid_filter_6_11(hash_out_valid_filter_6_11),
    .hash_out_6_12(hash_out_6_12),
    .hash_out_valid_filter_6_12(hash_out_valid_filter_6_12),
    .hash_out_6_13(hash_out_6_13),
    .hash_out_valid_filter_6_13(hash_out_valid_filter_6_13),
    .hash_out_6_14(hash_out_6_14),
    .hash_out_valid_filter_6_14(hash_out_valid_filter_6_14),
    .hash_out_6_15(hash_out_6_15),
    .hash_out_valid_filter_6_15(hash_out_valid_filter_6_15),
    .hash_out_6_16(hash_out_6_16),
    .hash_out_valid_filter_6_16(hash_out_valid_filter_6_16),
    .hash_out_6_17(hash_out_6_17),
    .hash_out_valid_filter_6_17(hash_out_valid_filter_6_17),
    .hash_out_6_18(hash_out_6_18),
    .hash_out_valid_filter_6_18(hash_out_valid_filter_6_18),
    .hash_out_6_19(hash_out_6_19),
    .hash_out_valid_filter_6_19(hash_out_valid_filter_6_19),
    .hash_out_6_20(hash_out_6_20),
    .hash_out_valid_filter_6_20(hash_out_valid_filter_6_20),
    .hash_out_6_21(hash_out_6_21),
    .hash_out_valid_filter_6_21(hash_out_valid_filter_6_21),
    .hash_out_6_22(hash_out_6_22),
    .hash_out_valid_filter_6_22(hash_out_valid_filter_6_22),
    .hash_out_6_23(hash_out_6_23),
    .hash_out_valid_filter_6_23(hash_out_valid_filter_6_23),
    .hash_out_6_24(hash_out_6_24),
    .hash_out_valid_filter_6_24(hash_out_valid_filter_6_24),
    .hash_out_6_25(hash_out_6_25),
    .hash_out_valid_filter_6_25(hash_out_valid_filter_6_25),
    .hash_out_6_26(hash_out_6_26),
    .hash_out_valid_filter_6_26(hash_out_valid_filter_6_26),
    .hash_out_6_27(hash_out_6_27),
    .hash_out_valid_filter_6_27(hash_out_valid_filter_6_27),
    .hash_out_6_28(hash_out_6_28),
    .hash_out_valid_filter_6_28(hash_out_valid_filter_6_28),
    .hash_out_6_29(hash_out_6_29),
    .hash_out_valid_filter_6_29(hash_out_valid_filter_6_29),
    .hash_out_6_30(hash_out_6_30),
    .hash_out_valid_filter_6_30(hash_out_valid_filter_6_30),
    .hash_out_6_31(hash_out_6_31),
    .hash_out_valid_filter_6_31(hash_out_valid_filter_6_31),
    .hash_out_7_0(hash_out_7_0),
    .hash_out_valid_filter_7_0(hash_out_valid_filter_7_0),
    .hash_out_7_1(hash_out_7_1),
    .hash_out_valid_filter_7_1(hash_out_valid_filter_7_1),
    .hash_out_7_2(hash_out_7_2),
    .hash_out_valid_filter_7_2(hash_out_valid_filter_7_2),
    .hash_out_7_3(hash_out_7_3),
    .hash_out_valid_filter_7_3(hash_out_valid_filter_7_3),
    .hash_out_7_4(hash_out_7_4),
    .hash_out_valid_filter_7_4(hash_out_valid_filter_7_4),
    .hash_out_7_5(hash_out_7_5),
    .hash_out_valid_filter_7_5(hash_out_valid_filter_7_5),
    .hash_out_7_6(hash_out_7_6),
    .hash_out_valid_filter_7_6(hash_out_valid_filter_7_6),
    .hash_out_7_7(hash_out_7_7),
    .hash_out_valid_filter_7_7(hash_out_valid_filter_7_7),
    .hash_out_7_8(hash_out_7_8),
    .hash_out_valid_filter_7_8(hash_out_valid_filter_7_8),
    .hash_out_7_9(hash_out_7_9),
    .hash_out_valid_filter_7_9(hash_out_valid_filter_7_9),
    .hash_out_7_10(hash_out_7_10),
    .hash_out_valid_filter_7_10(hash_out_valid_filter_7_10),
    .hash_out_7_11(hash_out_7_11),
    .hash_out_valid_filter_7_11(hash_out_valid_filter_7_11),
    .hash_out_7_12(hash_out_7_12),
    .hash_out_valid_filter_7_12(hash_out_valid_filter_7_12),
    .hash_out_7_13(hash_out_7_13),
    .hash_out_valid_filter_7_13(hash_out_valid_filter_7_13),
    .hash_out_7_14(hash_out_7_14),
    .hash_out_valid_filter_7_14(hash_out_valid_filter_7_14),
    .hash_out_7_15(hash_out_7_15),
    .hash_out_valid_filter_7_15(hash_out_valid_filter_7_15),
    .hash_out_7_16(hash_out_7_16),
    .hash_out_valid_filter_7_16(hash_out_valid_filter_7_16),
    .hash_out_7_17(hash_out_7_17),
    .hash_out_valid_filter_7_17(hash_out_valid_filter_7_17),
    .hash_out_7_18(hash_out_7_18),
    .hash_out_valid_filter_7_18(hash_out_valid_filter_7_18),
    .hash_out_7_19(hash_out_7_19),
    .hash_out_valid_filter_7_19(hash_out_valid_filter_7_19),
    .hash_out_7_20(hash_out_7_20),
    .hash_out_valid_filter_7_20(hash_out_valid_filter_7_20),
    .hash_out_7_21(hash_out_7_21),
    .hash_out_valid_filter_7_21(hash_out_valid_filter_7_21),
    .hash_out_7_22(hash_out_7_22),
    .hash_out_valid_filter_7_22(hash_out_valid_filter_7_22),
    .hash_out_7_23(hash_out_7_23),
    .hash_out_valid_filter_7_23(hash_out_valid_filter_7_23),
    .hash_out_7_24(hash_out_7_24),
    .hash_out_valid_filter_7_24(hash_out_valid_filter_7_24),
    .hash_out_7_25(hash_out_7_25),
    .hash_out_valid_filter_7_25(hash_out_valid_filter_7_25),
    .hash_out_7_26(hash_out_7_26),
    .hash_out_valid_filter_7_26(hash_out_valid_filter_7_26),
    .hash_out_7_27(hash_out_7_27),
    .hash_out_valid_filter_7_27(hash_out_valid_filter_7_27),
    .hash_out_7_28(hash_out_7_28),
    .hash_out_valid_filter_7_28(hash_out_valid_filter_7_28),
    .hash_out_7_29(hash_out_7_29),
    .hash_out_valid_filter_7_29(hash_out_valid_filter_7_29),
    .hash_out_7_30(hash_out_7_30),
    .hash_out_valid_filter_7_30(hash_out_valid_filter_7_30),
    .hash_out_7_31(hash_out_7_31),
    .hash_out_valid_filter_7_31(hash_out_valid_filter_7_31),
    .in_data(in_data_r2),
    .in_valid(in_valid_r2),
    .in_sop(in_sop_r2),
    .in_eop(in_eop_r2),
    .in_empty(in_empty_r2),
    .out_new_pkt(out_new_pkt)
);

//RuleID reduction logic
backend back(
    .clk(clk),
    .rst(rst),
    .din_0_0(din_0_0_r2),
    .din_valid_0_0(din_valid_0_0_r2),
    .din_almost_full_0_0(din_almost_full_0_0),
    .din_0_1(din_0_1_r2),
    .din_valid_0_1(din_valid_0_1_r2),
    .din_almost_full_0_1(din_almost_full_0_1),
    .din_0_2(din_0_2_r2),
    .din_valid_0_2(din_valid_0_2_r2),
    .din_almost_full_0_2(din_almost_full_0_2),
    .din_0_3(din_0_3_r2),
    .din_valid_0_3(din_valid_0_3_r2),
    .din_almost_full_0_3(din_almost_full_0_3),
    .din_0_4(din_0_4_r2),
    .din_valid_0_4(din_valid_0_4_r2),
    .din_almost_full_0_4(din_almost_full_0_4),
    .din_0_5(din_0_5_r2),
    .din_valid_0_5(din_valid_0_5_r2),
    .din_almost_full_0_5(din_almost_full_0_5),
    .din_0_6(din_0_6_r2),
    .din_valid_0_6(din_valid_0_6_r2),
    .din_almost_full_0_6(din_almost_full_0_6),
    .din_0_7(din_0_7_r2),
    .din_valid_0_7(din_valid_0_7_r2),
    .din_almost_full_0_7(din_almost_full_0_7),
    .din_0_8(din_0_8_r2),
    .din_valid_0_8(din_valid_0_8_r2),
    .din_almost_full_0_8(din_almost_full_0_8),
    .din_0_9(din_0_9_r2),
    .din_valid_0_9(din_valid_0_9_r2),
    .din_almost_full_0_9(din_almost_full_0_9),
    .din_0_10(din_0_10_r2),
    .din_valid_0_10(din_valid_0_10_r2),
    .din_almost_full_0_10(din_almost_full_0_10),
    .din_0_11(din_0_11_r2),
    .din_valid_0_11(din_valid_0_11_r2),
    .din_almost_full_0_11(din_almost_full_0_11),
    .din_0_12(din_0_12_r2),
    .din_valid_0_12(din_valid_0_12_r2),
    .din_almost_full_0_12(din_almost_full_0_12),
    .din_0_13(din_0_13_r2),
    .din_valid_0_13(din_valid_0_13_r2),
    .din_almost_full_0_13(din_almost_full_0_13),
    .din_0_14(din_0_14_r2),
    .din_valid_0_14(din_valid_0_14_r2),
    .din_almost_full_0_14(din_almost_full_0_14),
    .din_0_15(din_0_15_r2),
    .din_valid_0_15(din_valid_0_15_r2),
    .din_almost_full_0_15(din_almost_full_0_15),
    .din_0_16(din_0_16_r2),
    .din_valid_0_16(din_valid_0_16_r2),
    .din_almost_full_0_16(din_almost_full_0_16),
    .din_0_17(din_0_17_r2),
    .din_valid_0_17(din_valid_0_17_r2),
    .din_almost_full_0_17(din_almost_full_0_17),
    .din_0_18(din_0_18_r2),
    .din_valid_0_18(din_valid_0_18_r2),
    .din_almost_full_0_18(din_almost_full_0_18),
    .din_0_19(din_0_19_r2),
    .din_valid_0_19(din_valid_0_19_r2),
    .din_almost_full_0_19(din_almost_full_0_19),
    .din_0_20(din_0_20_r2),
    .din_valid_0_20(din_valid_0_20_r2),
    .din_almost_full_0_20(din_almost_full_0_20),
    .din_0_21(din_0_21_r2),
    .din_valid_0_21(din_valid_0_21_r2),
    .din_almost_full_0_21(din_almost_full_0_21),
    .din_0_22(din_0_22_r2),
    .din_valid_0_22(din_valid_0_22_r2),
    .din_almost_full_0_22(din_almost_full_0_22),
    .din_0_23(din_0_23_r2),
    .din_valid_0_23(din_valid_0_23_r2),
    .din_almost_full_0_23(din_almost_full_0_23),
    .din_0_24(din_0_24_r2),
    .din_valid_0_24(din_valid_0_24_r2),
    .din_almost_full_0_24(din_almost_full_0_24),
    .din_0_25(din_0_25_r2),
    .din_valid_0_25(din_valid_0_25_r2),
    .din_almost_full_0_25(din_almost_full_0_25),
    .din_0_26(din_0_26_r2),
    .din_valid_0_26(din_valid_0_26_r2),
    .din_almost_full_0_26(din_almost_full_0_26),
    .din_0_27(din_0_27_r2),
    .din_valid_0_27(din_valid_0_27_r2),
    .din_almost_full_0_27(din_almost_full_0_27),
    .din_0_28(din_0_28_r2),
    .din_valid_0_28(din_valid_0_28_r2),
    .din_almost_full_0_28(din_almost_full_0_28),
    .din_0_29(din_0_29_r2),
    .din_valid_0_29(din_valid_0_29_r2),
    .din_almost_full_0_29(din_almost_full_0_29),
    .din_0_30(din_0_30_r2),
    .din_valid_0_30(din_valid_0_30_r2),
    .din_almost_full_0_30(din_almost_full_0_30),
    .din_0_31(din_0_31_r2),
    .din_valid_0_31(din_valid_0_31_r2),
    .din_almost_full_0_31(din_almost_full_0_31),
    .din_1_0(din_1_0_r2),
    .din_valid_1_0(din_valid_1_0_r2),
    .din_almost_full_1_0(din_almost_full_1_0),
    .din_1_1(din_1_1_r2),
    .din_valid_1_1(din_valid_1_1_r2),
    .din_almost_full_1_1(din_almost_full_1_1),
    .din_1_2(din_1_2_r2),
    .din_valid_1_2(din_valid_1_2_r2),
    .din_almost_full_1_2(din_almost_full_1_2),
    .din_1_3(din_1_3_r2),
    .din_valid_1_3(din_valid_1_3_r2),
    .din_almost_full_1_3(din_almost_full_1_3),
    .din_1_4(din_1_4_r2),
    .din_valid_1_4(din_valid_1_4_r2),
    .din_almost_full_1_4(din_almost_full_1_4),
    .din_1_5(din_1_5_r2),
    .din_valid_1_5(din_valid_1_5_r2),
    .din_almost_full_1_5(din_almost_full_1_5),
    .din_1_6(din_1_6_r2),
    .din_valid_1_6(din_valid_1_6_r2),
    .din_almost_full_1_6(din_almost_full_1_6),
    .din_1_7(din_1_7_r2),
    .din_valid_1_7(din_valid_1_7_r2),
    .din_almost_full_1_7(din_almost_full_1_7),
    .din_1_8(din_1_8_r2),
    .din_valid_1_8(din_valid_1_8_r2),
    .din_almost_full_1_8(din_almost_full_1_8),
    .din_1_9(din_1_9_r2),
    .din_valid_1_9(din_valid_1_9_r2),
    .din_almost_full_1_9(din_almost_full_1_9),
    .din_1_10(din_1_10_r2),
    .din_valid_1_10(din_valid_1_10_r2),
    .din_almost_full_1_10(din_almost_full_1_10),
    .din_1_11(din_1_11_r2),
    .din_valid_1_11(din_valid_1_11_r2),
    .din_almost_full_1_11(din_almost_full_1_11),
    .din_1_12(din_1_12_r2),
    .din_valid_1_12(din_valid_1_12_r2),
    .din_almost_full_1_12(din_almost_full_1_12),
    .din_1_13(din_1_13_r2),
    .din_valid_1_13(din_valid_1_13_r2),
    .din_almost_full_1_13(din_almost_full_1_13),
    .din_1_14(din_1_14_r2),
    .din_valid_1_14(din_valid_1_14_r2),
    .din_almost_full_1_14(din_almost_full_1_14),
    .din_1_15(din_1_15_r2),
    .din_valid_1_15(din_valid_1_15_r2),
    .din_almost_full_1_15(din_almost_full_1_15),
    .din_1_16(din_1_16_r2),
    .din_valid_1_16(din_valid_1_16_r2),
    .din_almost_full_1_16(din_almost_full_1_16),
    .din_1_17(din_1_17_r2),
    .din_valid_1_17(din_valid_1_17_r2),
    .din_almost_full_1_17(din_almost_full_1_17),
    .din_1_18(din_1_18_r2),
    .din_valid_1_18(din_valid_1_18_r2),
    .din_almost_full_1_18(din_almost_full_1_18),
    .din_1_19(din_1_19_r2),
    .din_valid_1_19(din_valid_1_19_r2),
    .din_almost_full_1_19(din_almost_full_1_19),
    .din_1_20(din_1_20_r2),
    .din_valid_1_20(din_valid_1_20_r2),
    .din_almost_full_1_20(din_almost_full_1_20),
    .din_1_21(din_1_21_r2),
    .din_valid_1_21(din_valid_1_21_r2),
    .din_almost_full_1_21(din_almost_full_1_21),
    .din_1_22(din_1_22_r2),
    .din_valid_1_22(din_valid_1_22_r2),
    .din_almost_full_1_22(din_almost_full_1_22),
    .din_1_23(din_1_23_r2),
    .din_valid_1_23(din_valid_1_23_r2),
    .din_almost_full_1_23(din_almost_full_1_23),
    .din_1_24(din_1_24_r2),
    .din_valid_1_24(din_valid_1_24_r2),
    .din_almost_full_1_24(din_almost_full_1_24),
    .din_1_25(din_1_25_r2),
    .din_valid_1_25(din_valid_1_25_r2),
    .din_almost_full_1_25(din_almost_full_1_25),
    .din_1_26(din_1_26_r2),
    .din_valid_1_26(din_valid_1_26_r2),
    .din_almost_full_1_26(din_almost_full_1_26),
    .din_1_27(din_1_27_r2),
    .din_valid_1_27(din_valid_1_27_r2),
    .din_almost_full_1_27(din_almost_full_1_27),
    .din_1_28(din_1_28_r2),
    .din_valid_1_28(din_valid_1_28_r2),
    .din_almost_full_1_28(din_almost_full_1_28),
    .din_1_29(din_1_29_r2),
    .din_valid_1_29(din_valid_1_29_r2),
    .din_almost_full_1_29(din_almost_full_1_29),
    .din_1_30(din_1_30_r2),
    .din_valid_1_30(din_valid_1_30_r2),
    .din_almost_full_1_30(din_almost_full_1_30),
    .din_1_31(din_1_31_r2),
    .din_valid_1_31(din_valid_1_31_r2),
    .din_almost_full_1_31(din_almost_full_1_31),
    .din_2_0(din_2_0_r2),
    .din_valid_2_0(din_valid_2_0_r2),
    .din_almost_full_2_0(din_almost_full_2_0),
    .din_2_1(din_2_1_r2),
    .din_valid_2_1(din_valid_2_1_r2),
    .din_almost_full_2_1(din_almost_full_2_1),
    .din_2_2(din_2_2_r2),
    .din_valid_2_2(din_valid_2_2_r2),
    .din_almost_full_2_2(din_almost_full_2_2),
    .din_2_3(din_2_3_r2),
    .din_valid_2_3(din_valid_2_3_r2),
    .din_almost_full_2_3(din_almost_full_2_3),
    .din_2_4(din_2_4_r2),
    .din_valid_2_4(din_valid_2_4_r2),
    .din_almost_full_2_4(din_almost_full_2_4),
    .din_2_5(din_2_5_r2),
    .din_valid_2_5(din_valid_2_5_r2),
    .din_almost_full_2_5(din_almost_full_2_5),
    .din_2_6(din_2_6_r2),
    .din_valid_2_6(din_valid_2_6_r2),
    .din_almost_full_2_6(din_almost_full_2_6),
    .din_2_7(din_2_7_r2),
    .din_valid_2_7(din_valid_2_7_r2),
    .din_almost_full_2_7(din_almost_full_2_7),
    .din_2_8(din_2_8_r2),
    .din_valid_2_8(din_valid_2_8_r2),
    .din_almost_full_2_8(din_almost_full_2_8),
    .din_2_9(din_2_9_r2),
    .din_valid_2_9(din_valid_2_9_r2),
    .din_almost_full_2_9(din_almost_full_2_9),
    .din_2_10(din_2_10_r2),
    .din_valid_2_10(din_valid_2_10_r2),
    .din_almost_full_2_10(din_almost_full_2_10),
    .din_2_11(din_2_11_r2),
    .din_valid_2_11(din_valid_2_11_r2),
    .din_almost_full_2_11(din_almost_full_2_11),
    .din_2_12(din_2_12_r2),
    .din_valid_2_12(din_valid_2_12_r2),
    .din_almost_full_2_12(din_almost_full_2_12),
    .din_2_13(din_2_13_r2),
    .din_valid_2_13(din_valid_2_13_r2),
    .din_almost_full_2_13(din_almost_full_2_13),
    .din_2_14(din_2_14_r2),
    .din_valid_2_14(din_valid_2_14_r2),
    .din_almost_full_2_14(din_almost_full_2_14),
    .din_2_15(din_2_15_r2),
    .din_valid_2_15(din_valid_2_15_r2),
    .din_almost_full_2_15(din_almost_full_2_15),
    .din_2_16(din_2_16_r2),
    .din_valid_2_16(din_valid_2_16_r2),
    .din_almost_full_2_16(din_almost_full_2_16),
    .din_2_17(din_2_17_r2),
    .din_valid_2_17(din_valid_2_17_r2),
    .din_almost_full_2_17(din_almost_full_2_17),
    .din_2_18(din_2_18_r2),
    .din_valid_2_18(din_valid_2_18_r2),
    .din_almost_full_2_18(din_almost_full_2_18),
    .din_2_19(din_2_19_r2),
    .din_valid_2_19(din_valid_2_19_r2),
    .din_almost_full_2_19(din_almost_full_2_19),
    .din_2_20(din_2_20_r2),
    .din_valid_2_20(din_valid_2_20_r2),
    .din_almost_full_2_20(din_almost_full_2_20),
    .din_2_21(din_2_21_r2),
    .din_valid_2_21(din_valid_2_21_r2),
    .din_almost_full_2_21(din_almost_full_2_21),
    .din_2_22(din_2_22_r2),
    .din_valid_2_22(din_valid_2_22_r2),
    .din_almost_full_2_22(din_almost_full_2_22),
    .din_2_23(din_2_23_r2),
    .din_valid_2_23(din_valid_2_23_r2),
    .din_almost_full_2_23(din_almost_full_2_23),
    .din_2_24(din_2_24_r2),
    .din_valid_2_24(din_valid_2_24_r2),
    .din_almost_full_2_24(din_almost_full_2_24),
    .din_2_25(din_2_25_r2),
    .din_valid_2_25(din_valid_2_25_r2),
    .din_almost_full_2_25(din_almost_full_2_25),
    .din_2_26(din_2_26_r2),
    .din_valid_2_26(din_valid_2_26_r2),
    .din_almost_full_2_26(din_almost_full_2_26),
    .din_2_27(din_2_27_r2),
    .din_valid_2_27(din_valid_2_27_r2),
    .din_almost_full_2_27(din_almost_full_2_27),
    .din_2_28(din_2_28_r2),
    .din_valid_2_28(din_valid_2_28_r2),
    .din_almost_full_2_28(din_almost_full_2_28),
    .din_2_29(din_2_29_r2),
    .din_valid_2_29(din_valid_2_29_r2),
    .din_almost_full_2_29(din_almost_full_2_29),
    .din_2_30(din_2_30_r2),
    .din_valid_2_30(din_valid_2_30_r2),
    .din_almost_full_2_30(din_almost_full_2_30),
    .din_2_31(din_2_31_r2),
    .din_valid_2_31(din_valid_2_31_r2),
    .din_almost_full_2_31(din_almost_full_2_31),
    .din_3_0(din_3_0_r2),
    .din_valid_3_0(din_valid_3_0_r2),
    .din_almost_full_3_0(din_almost_full_3_0),
    .din_3_1(din_3_1_r2),
    .din_valid_3_1(din_valid_3_1_r2),
    .din_almost_full_3_1(din_almost_full_3_1),
    .din_3_2(din_3_2_r2),
    .din_valid_3_2(din_valid_3_2_r2),
    .din_almost_full_3_2(din_almost_full_3_2),
    .din_3_3(din_3_3_r2),
    .din_valid_3_3(din_valid_3_3_r2),
    .din_almost_full_3_3(din_almost_full_3_3),
    .din_3_4(din_3_4_r2),
    .din_valid_3_4(din_valid_3_4_r2),
    .din_almost_full_3_4(din_almost_full_3_4),
    .din_3_5(din_3_5_r2),
    .din_valid_3_5(din_valid_3_5_r2),
    .din_almost_full_3_5(din_almost_full_3_5),
    .din_3_6(din_3_6_r2),
    .din_valid_3_6(din_valid_3_6_r2),
    .din_almost_full_3_6(din_almost_full_3_6),
    .din_3_7(din_3_7_r2),
    .din_valid_3_7(din_valid_3_7_r2),
    .din_almost_full_3_7(din_almost_full_3_7),
    .din_3_8(din_3_8_r2),
    .din_valid_3_8(din_valid_3_8_r2),
    .din_almost_full_3_8(din_almost_full_3_8),
    .din_3_9(din_3_9_r2),
    .din_valid_3_9(din_valid_3_9_r2),
    .din_almost_full_3_9(din_almost_full_3_9),
    .din_3_10(din_3_10_r2),
    .din_valid_3_10(din_valid_3_10_r2),
    .din_almost_full_3_10(din_almost_full_3_10),
    .din_3_11(din_3_11_r2),
    .din_valid_3_11(din_valid_3_11_r2),
    .din_almost_full_3_11(din_almost_full_3_11),
    .din_3_12(din_3_12_r2),
    .din_valid_3_12(din_valid_3_12_r2),
    .din_almost_full_3_12(din_almost_full_3_12),
    .din_3_13(din_3_13_r2),
    .din_valid_3_13(din_valid_3_13_r2),
    .din_almost_full_3_13(din_almost_full_3_13),
    .din_3_14(din_3_14_r2),
    .din_valid_3_14(din_valid_3_14_r2),
    .din_almost_full_3_14(din_almost_full_3_14),
    .din_3_15(din_3_15_r2),
    .din_valid_3_15(din_valid_3_15_r2),
    .din_almost_full_3_15(din_almost_full_3_15),
    .din_3_16(din_3_16_r2),
    .din_valid_3_16(din_valid_3_16_r2),
    .din_almost_full_3_16(din_almost_full_3_16),
    .din_3_17(din_3_17_r2),
    .din_valid_3_17(din_valid_3_17_r2),
    .din_almost_full_3_17(din_almost_full_3_17),
    .din_3_18(din_3_18_r2),
    .din_valid_3_18(din_valid_3_18_r2),
    .din_almost_full_3_18(din_almost_full_3_18),
    .din_3_19(din_3_19_r2),
    .din_valid_3_19(din_valid_3_19_r2),
    .din_almost_full_3_19(din_almost_full_3_19),
    .din_3_20(din_3_20_r2),
    .din_valid_3_20(din_valid_3_20_r2),
    .din_almost_full_3_20(din_almost_full_3_20),
    .din_3_21(din_3_21_r2),
    .din_valid_3_21(din_valid_3_21_r2),
    .din_almost_full_3_21(din_almost_full_3_21),
    .din_3_22(din_3_22_r2),
    .din_valid_3_22(din_valid_3_22_r2),
    .din_almost_full_3_22(din_almost_full_3_22),
    .din_3_23(din_3_23_r2),
    .din_valid_3_23(din_valid_3_23_r2),
    .din_almost_full_3_23(din_almost_full_3_23),
    .din_3_24(din_3_24_r2),
    .din_valid_3_24(din_valid_3_24_r2),
    .din_almost_full_3_24(din_almost_full_3_24),
    .din_3_25(din_3_25_r2),
    .din_valid_3_25(din_valid_3_25_r2),
    .din_almost_full_3_25(din_almost_full_3_25),
    .din_3_26(din_3_26_r2),
    .din_valid_3_26(din_valid_3_26_r2),
    .din_almost_full_3_26(din_almost_full_3_26),
    .din_3_27(din_3_27_r2),
    .din_valid_3_27(din_valid_3_27_r2),
    .din_almost_full_3_27(din_almost_full_3_27),
    .din_3_28(din_3_28_r2),
    .din_valid_3_28(din_valid_3_28_r2),
    .din_almost_full_3_28(din_almost_full_3_28),
    .din_3_29(din_3_29_r2),
    .din_valid_3_29(din_valid_3_29_r2),
    .din_almost_full_3_29(din_almost_full_3_29),
    .din_3_30(din_3_30_r2),
    .din_valid_3_30(din_valid_3_30_r2),
    .din_almost_full_3_30(din_almost_full_3_30),
    .din_3_31(din_3_31_r2),
    .din_valid_3_31(din_valid_3_31_r2),
    .din_almost_full_3_31(din_almost_full_3_31),
    .din_4_0(din_4_0_r2),
    .din_valid_4_0(din_valid_4_0_r2),
    .din_almost_full_4_0(din_almost_full_4_0),
    .din_4_1(din_4_1_r2),
    .din_valid_4_1(din_valid_4_1_r2),
    .din_almost_full_4_1(din_almost_full_4_1),
    .din_4_2(din_4_2_r2),
    .din_valid_4_2(din_valid_4_2_r2),
    .din_almost_full_4_2(din_almost_full_4_2),
    .din_4_3(din_4_3_r2),
    .din_valid_4_3(din_valid_4_3_r2),
    .din_almost_full_4_3(din_almost_full_4_3),
    .din_4_4(din_4_4_r2),
    .din_valid_4_4(din_valid_4_4_r2),
    .din_almost_full_4_4(din_almost_full_4_4),
    .din_4_5(din_4_5_r2),
    .din_valid_4_5(din_valid_4_5_r2),
    .din_almost_full_4_5(din_almost_full_4_5),
    .din_4_6(din_4_6_r2),
    .din_valid_4_6(din_valid_4_6_r2),
    .din_almost_full_4_6(din_almost_full_4_6),
    .din_4_7(din_4_7_r2),
    .din_valid_4_7(din_valid_4_7_r2),
    .din_almost_full_4_7(din_almost_full_4_7),
    .din_4_8(din_4_8_r2),
    .din_valid_4_8(din_valid_4_8_r2),
    .din_almost_full_4_8(din_almost_full_4_8),
    .din_4_9(din_4_9_r2),
    .din_valid_4_9(din_valid_4_9_r2),
    .din_almost_full_4_9(din_almost_full_4_9),
    .din_4_10(din_4_10_r2),
    .din_valid_4_10(din_valid_4_10_r2),
    .din_almost_full_4_10(din_almost_full_4_10),
    .din_4_11(din_4_11_r2),
    .din_valid_4_11(din_valid_4_11_r2),
    .din_almost_full_4_11(din_almost_full_4_11),
    .din_4_12(din_4_12_r2),
    .din_valid_4_12(din_valid_4_12_r2),
    .din_almost_full_4_12(din_almost_full_4_12),
    .din_4_13(din_4_13_r2),
    .din_valid_4_13(din_valid_4_13_r2),
    .din_almost_full_4_13(din_almost_full_4_13),
    .din_4_14(din_4_14_r2),
    .din_valid_4_14(din_valid_4_14_r2),
    .din_almost_full_4_14(din_almost_full_4_14),
    .din_4_15(din_4_15_r2),
    .din_valid_4_15(din_valid_4_15_r2),
    .din_almost_full_4_15(din_almost_full_4_15),
    .din_4_16(din_4_16_r2),
    .din_valid_4_16(din_valid_4_16_r2),
    .din_almost_full_4_16(din_almost_full_4_16),
    .din_4_17(din_4_17_r2),
    .din_valid_4_17(din_valid_4_17_r2),
    .din_almost_full_4_17(din_almost_full_4_17),
    .din_4_18(din_4_18_r2),
    .din_valid_4_18(din_valid_4_18_r2),
    .din_almost_full_4_18(din_almost_full_4_18),
    .din_4_19(din_4_19_r2),
    .din_valid_4_19(din_valid_4_19_r2),
    .din_almost_full_4_19(din_almost_full_4_19),
    .din_4_20(din_4_20_r2),
    .din_valid_4_20(din_valid_4_20_r2),
    .din_almost_full_4_20(din_almost_full_4_20),
    .din_4_21(din_4_21_r2),
    .din_valid_4_21(din_valid_4_21_r2),
    .din_almost_full_4_21(din_almost_full_4_21),
    .din_4_22(din_4_22_r2),
    .din_valid_4_22(din_valid_4_22_r2),
    .din_almost_full_4_22(din_almost_full_4_22),
    .din_4_23(din_4_23_r2),
    .din_valid_4_23(din_valid_4_23_r2),
    .din_almost_full_4_23(din_almost_full_4_23),
    .din_4_24(din_4_24_r2),
    .din_valid_4_24(din_valid_4_24_r2),
    .din_almost_full_4_24(din_almost_full_4_24),
    .din_4_25(din_4_25_r2),
    .din_valid_4_25(din_valid_4_25_r2),
    .din_almost_full_4_25(din_almost_full_4_25),
    .din_4_26(din_4_26_r2),
    .din_valid_4_26(din_valid_4_26_r2),
    .din_almost_full_4_26(din_almost_full_4_26),
    .din_4_27(din_4_27_r2),
    .din_valid_4_27(din_valid_4_27_r2),
    .din_almost_full_4_27(din_almost_full_4_27),
    .din_4_28(din_4_28_r2),
    .din_valid_4_28(din_valid_4_28_r2),
    .din_almost_full_4_28(din_almost_full_4_28),
    .din_4_29(din_4_29_r2),
    .din_valid_4_29(din_valid_4_29_r2),
    .din_almost_full_4_29(din_almost_full_4_29),
    .din_4_30(din_4_30_r2),
    .din_valid_4_30(din_valid_4_30_r2),
    .din_almost_full_4_30(din_almost_full_4_30),
    .din_4_31(din_4_31_r2),
    .din_valid_4_31(din_valid_4_31_r2),
    .din_almost_full_4_31(din_almost_full_4_31),
    .din_5_0(din_5_0_r2),
    .din_valid_5_0(din_valid_5_0_r2),
    .din_almost_full_5_0(din_almost_full_5_0),
    .din_5_1(din_5_1_r2),
    .din_valid_5_1(din_valid_5_1_r2),
    .din_almost_full_5_1(din_almost_full_5_1),
    .din_5_2(din_5_2_r2),
    .din_valid_5_2(din_valid_5_2_r2),
    .din_almost_full_5_2(din_almost_full_5_2),
    .din_5_3(din_5_3_r2),
    .din_valid_5_3(din_valid_5_3_r2),
    .din_almost_full_5_3(din_almost_full_5_3),
    .din_5_4(din_5_4_r2),
    .din_valid_5_4(din_valid_5_4_r2),
    .din_almost_full_5_4(din_almost_full_5_4),
    .din_5_5(din_5_5_r2),
    .din_valid_5_5(din_valid_5_5_r2),
    .din_almost_full_5_5(din_almost_full_5_5),
    .din_5_6(din_5_6_r2),
    .din_valid_5_6(din_valid_5_6_r2),
    .din_almost_full_5_6(din_almost_full_5_6),
    .din_5_7(din_5_7_r2),
    .din_valid_5_7(din_valid_5_7_r2),
    .din_almost_full_5_7(din_almost_full_5_7),
    .din_5_8(din_5_8_r2),
    .din_valid_5_8(din_valid_5_8_r2),
    .din_almost_full_5_8(din_almost_full_5_8),
    .din_5_9(din_5_9_r2),
    .din_valid_5_9(din_valid_5_9_r2),
    .din_almost_full_5_9(din_almost_full_5_9),
    .din_5_10(din_5_10_r2),
    .din_valid_5_10(din_valid_5_10_r2),
    .din_almost_full_5_10(din_almost_full_5_10),
    .din_5_11(din_5_11_r2),
    .din_valid_5_11(din_valid_5_11_r2),
    .din_almost_full_5_11(din_almost_full_5_11),
    .din_5_12(din_5_12_r2),
    .din_valid_5_12(din_valid_5_12_r2),
    .din_almost_full_5_12(din_almost_full_5_12),
    .din_5_13(din_5_13_r2),
    .din_valid_5_13(din_valid_5_13_r2),
    .din_almost_full_5_13(din_almost_full_5_13),
    .din_5_14(din_5_14_r2),
    .din_valid_5_14(din_valid_5_14_r2),
    .din_almost_full_5_14(din_almost_full_5_14),
    .din_5_15(din_5_15_r2),
    .din_valid_5_15(din_valid_5_15_r2),
    .din_almost_full_5_15(din_almost_full_5_15),
    .din_5_16(din_5_16_r2),
    .din_valid_5_16(din_valid_5_16_r2),
    .din_almost_full_5_16(din_almost_full_5_16),
    .din_5_17(din_5_17_r2),
    .din_valid_5_17(din_valid_5_17_r2),
    .din_almost_full_5_17(din_almost_full_5_17),
    .din_5_18(din_5_18_r2),
    .din_valid_5_18(din_valid_5_18_r2),
    .din_almost_full_5_18(din_almost_full_5_18),
    .din_5_19(din_5_19_r2),
    .din_valid_5_19(din_valid_5_19_r2),
    .din_almost_full_5_19(din_almost_full_5_19),
    .din_5_20(din_5_20_r2),
    .din_valid_5_20(din_valid_5_20_r2),
    .din_almost_full_5_20(din_almost_full_5_20),
    .din_5_21(din_5_21_r2),
    .din_valid_5_21(din_valid_5_21_r2),
    .din_almost_full_5_21(din_almost_full_5_21),
    .din_5_22(din_5_22_r2),
    .din_valid_5_22(din_valid_5_22_r2),
    .din_almost_full_5_22(din_almost_full_5_22),
    .din_5_23(din_5_23_r2),
    .din_valid_5_23(din_valid_5_23_r2),
    .din_almost_full_5_23(din_almost_full_5_23),
    .din_5_24(din_5_24_r2),
    .din_valid_5_24(din_valid_5_24_r2),
    .din_almost_full_5_24(din_almost_full_5_24),
    .din_5_25(din_5_25_r2),
    .din_valid_5_25(din_valid_5_25_r2),
    .din_almost_full_5_25(din_almost_full_5_25),
    .din_5_26(din_5_26_r2),
    .din_valid_5_26(din_valid_5_26_r2),
    .din_almost_full_5_26(din_almost_full_5_26),
    .din_5_27(din_5_27_r2),
    .din_valid_5_27(din_valid_5_27_r2),
    .din_almost_full_5_27(din_almost_full_5_27),
    .din_5_28(din_5_28_r2),
    .din_valid_5_28(din_valid_5_28_r2),
    .din_almost_full_5_28(din_almost_full_5_28),
    .din_5_29(din_5_29_r2),
    .din_valid_5_29(din_valid_5_29_r2),
    .din_almost_full_5_29(din_almost_full_5_29),
    .din_5_30(din_5_30_r2),
    .din_valid_5_30(din_valid_5_30_r2),
    .din_almost_full_5_30(din_almost_full_5_30),
    .din_5_31(din_5_31_r2),
    .din_valid_5_31(din_valid_5_31_r2),
    .din_almost_full_5_31(din_almost_full_5_31),
    .din_6_0(din_6_0_r2),
    .din_valid_6_0(din_valid_6_0_r2),
    .din_almost_full_6_0(din_almost_full_6_0),
    .din_6_1(din_6_1_r2),
    .din_valid_6_1(din_valid_6_1_r2),
    .din_almost_full_6_1(din_almost_full_6_1),
    .din_6_2(din_6_2_r2),
    .din_valid_6_2(din_valid_6_2_r2),
    .din_almost_full_6_2(din_almost_full_6_2),
    .din_6_3(din_6_3_r2),
    .din_valid_6_3(din_valid_6_3_r2),
    .din_almost_full_6_3(din_almost_full_6_3),
    .din_6_4(din_6_4_r2),
    .din_valid_6_4(din_valid_6_4_r2),
    .din_almost_full_6_4(din_almost_full_6_4),
    .din_6_5(din_6_5_r2),
    .din_valid_6_5(din_valid_6_5_r2),
    .din_almost_full_6_5(din_almost_full_6_5),
    .din_6_6(din_6_6_r2),
    .din_valid_6_6(din_valid_6_6_r2),
    .din_almost_full_6_6(din_almost_full_6_6),
    .din_6_7(din_6_7_r2),
    .din_valid_6_7(din_valid_6_7_r2),
    .din_almost_full_6_7(din_almost_full_6_7),
    .din_6_8(din_6_8_r2),
    .din_valid_6_8(din_valid_6_8_r2),
    .din_almost_full_6_8(din_almost_full_6_8),
    .din_6_9(din_6_9_r2),
    .din_valid_6_9(din_valid_6_9_r2),
    .din_almost_full_6_9(din_almost_full_6_9),
    .din_6_10(din_6_10_r2),
    .din_valid_6_10(din_valid_6_10_r2),
    .din_almost_full_6_10(din_almost_full_6_10),
    .din_6_11(din_6_11_r2),
    .din_valid_6_11(din_valid_6_11_r2),
    .din_almost_full_6_11(din_almost_full_6_11),
    .din_6_12(din_6_12_r2),
    .din_valid_6_12(din_valid_6_12_r2),
    .din_almost_full_6_12(din_almost_full_6_12),
    .din_6_13(din_6_13_r2),
    .din_valid_6_13(din_valid_6_13_r2),
    .din_almost_full_6_13(din_almost_full_6_13),
    .din_6_14(din_6_14_r2),
    .din_valid_6_14(din_valid_6_14_r2),
    .din_almost_full_6_14(din_almost_full_6_14),
    .din_6_15(din_6_15_r2),
    .din_valid_6_15(din_valid_6_15_r2),
    .din_almost_full_6_15(din_almost_full_6_15),
    .din_6_16(din_6_16_r2),
    .din_valid_6_16(din_valid_6_16_r2),
    .din_almost_full_6_16(din_almost_full_6_16),
    .din_6_17(din_6_17_r2),
    .din_valid_6_17(din_valid_6_17_r2),
    .din_almost_full_6_17(din_almost_full_6_17),
    .din_6_18(din_6_18_r2),
    .din_valid_6_18(din_valid_6_18_r2),
    .din_almost_full_6_18(din_almost_full_6_18),
    .din_6_19(din_6_19_r2),
    .din_valid_6_19(din_valid_6_19_r2),
    .din_almost_full_6_19(din_almost_full_6_19),
    .din_6_20(din_6_20_r2),
    .din_valid_6_20(din_valid_6_20_r2),
    .din_almost_full_6_20(din_almost_full_6_20),
    .din_6_21(din_6_21_r2),
    .din_valid_6_21(din_valid_6_21_r2),
    .din_almost_full_6_21(din_almost_full_6_21),
    .din_6_22(din_6_22_r2),
    .din_valid_6_22(din_valid_6_22_r2),
    .din_almost_full_6_22(din_almost_full_6_22),
    .din_6_23(din_6_23_r2),
    .din_valid_6_23(din_valid_6_23_r2),
    .din_almost_full_6_23(din_almost_full_6_23),
    .din_6_24(din_6_24_r2),
    .din_valid_6_24(din_valid_6_24_r2),
    .din_almost_full_6_24(din_almost_full_6_24),
    .din_6_25(din_6_25_r2),
    .din_valid_6_25(din_valid_6_25_r2),
    .din_almost_full_6_25(din_almost_full_6_25),
    .din_6_26(din_6_26_r2),
    .din_valid_6_26(din_valid_6_26_r2),
    .din_almost_full_6_26(din_almost_full_6_26),
    .din_6_27(din_6_27_r2),
    .din_valid_6_27(din_valid_6_27_r2),
    .din_almost_full_6_27(din_almost_full_6_27),
    .din_6_28(din_6_28_r2),
    .din_valid_6_28(din_valid_6_28_r2),
    .din_almost_full_6_28(din_almost_full_6_28),
    .din_6_29(din_6_29_r2),
    .din_valid_6_29(din_valid_6_29_r2),
    .din_almost_full_6_29(din_almost_full_6_29),
    .din_6_30(din_6_30_r2),
    .din_valid_6_30(din_valid_6_30_r2),
    .din_almost_full_6_30(din_almost_full_6_30),
    .din_6_31(din_6_31_r2),
    .din_valid_6_31(din_valid_6_31_r2),
    .din_almost_full_6_31(din_almost_full_6_31),
    .din_7_0(din_7_0_r2),
    .din_valid_7_0(din_valid_7_0_r2),
    .din_almost_full_7_0(din_almost_full_7_0),
    .din_7_1(din_7_1_r2),
    .din_valid_7_1(din_valid_7_1_r2),
    .din_almost_full_7_1(din_almost_full_7_1),
    .din_7_2(din_7_2_r2),
    .din_valid_7_2(din_valid_7_2_r2),
    .din_almost_full_7_2(din_almost_full_7_2),
    .din_7_3(din_7_3_r2),
    .din_valid_7_3(din_valid_7_3_r2),
    .din_almost_full_7_3(din_almost_full_7_3),
    .din_7_4(din_7_4_r2),
    .din_valid_7_4(din_valid_7_4_r2),
    .din_almost_full_7_4(din_almost_full_7_4),
    .din_7_5(din_7_5_r2),
    .din_valid_7_5(din_valid_7_5_r2),
    .din_almost_full_7_5(din_almost_full_7_5),
    .din_7_6(din_7_6_r2),
    .din_valid_7_6(din_valid_7_6_r2),
    .din_almost_full_7_6(din_almost_full_7_6),
    .din_7_7(din_7_7_r2),
    .din_valid_7_7(din_valid_7_7_r2),
    .din_almost_full_7_7(din_almost_full_7_7),
    .din_7_8(din_7_8_r2),
    .din_valid_7_8(din_valid_7_8_r2),
    .din_almost_full_7_8(din_almost_full_7_8),
    .din_7_9(din_7_9_r2),
    .din_valid_7_9(din_valid_7_9_r2),
    .din_almost_full_7_9(din_almost_full_7_9),
    .din_7_10(din_7_10_r2),
    .din_valid_7_10(din_valid_7_10_r2),
    .din_almost_full_7_10(din_almost_full_7_10),
    .din_7_11(din_7_11_r2),
    .din_valid_7_11(din_valid_7_11_r2),
    .din_almost_full_7_11(din_almost_full_7_11),
    .din_7_12(din_7_12_r2),
    .din_valid_7_12(din_valid_7_12_r2),
    .din_almost_full_7_12(din_almost_full_7_12),
    .din_7_13(din_7_13_r2),
    .din_valid_7_13(din_valid_7_13_r2),
    .din_almost_full_7_13(din_almost_full_7_13),
    .din_7_14(din_7_14_r2),
    .din_valid_7_14(din_valid_7_14_r2),
    .din_almost_full_7_14(din_almost_full_7_14),
    .din_7_15(din_7_15_r2),
    .din_valid_7_15(din_valid_7_15_r2),
    .din_almost_full_7_15(din_almost_full_7_15),
    .din_7_16(din_7_16_r2),
    .din_valid_7_16(din_valid_7_16_r2),
    .din_almost_full_7_16(din_almost_full_7_16),
    .din_7_17(din_7_17_r2),
    .din_valid_7_17(din_valid_7_17_r2),
    .din_almost_full_7_17(din_almost_full_7_17),
    .din_7_18(din_7_18_r2),
    .din_valid_7_18(din_valid_7_18_r2),
    .din_almost_full_7_18(din_almost_full_7_18),
    .din_7_19(din_7_19_r2),
    .din_valid_7_19(din_valid_7_19_r2),
    .din_almost_full_7_19(din_almost_full_7_19),
    .din_7_20(din_7_20_r2),
    .din_valid_7_20(din_valid_7_20_r2),
    .din_almost_full_7_20(din_almost_full_7_20),
    .din_7_21(din_7_21_r2),
    .din_valid_7_21(din_valid_7_21_r2),
    .din_almost_full_7_21(din_almost_full_7_21),
    .din_7_22(din_7_22_r2),
    .din_valid_7_22(din_valid_7_22_r2),
    .din_almost_full_7_22(din_almost_full_7_22),
    .din_7_23(din_7_23_r2),
    .din_valid_7_23(din_valid_7_23_r2),
    .din_almost_full_7_23(din_almost_full_7_23),
    .din_7_24(din_7_24_r2),
    .din_valid_7_24(din_valid_7_24_r2),
    .din_almost_full_7_24(din_almost_full_7_24),
    .din_7_25(din_7_25_r2),
    .din_valid_7_25(din_valid_7_25_r2),
    .din_almost_full_7_25(din_almost_full_7_25),
    .din_7_26(din_7_26_r2),
    .din_valid_7_26(din_valid_7_26_r2),
    .din_almost_full_7_26(din_almost_full_7_26),
    .din_7_27(din_7_27_r2),
    .din_valid_7_27(din_valid_7_27_r2),
    .din_almost_full_7_27(din_almost_full_7_27),
    .din_7_28(din_7_28_r2),
    .din_valid_7_28(din_valid_7_28_r2),
    .din_almost_full_7_28(din_almost_full_7_28),
    .din_7_29(din_7_29_r2),
    .din_valid_7_29(din_valid_7_29_r2),
    .din_almost_full_7_29(din_almost_full_7_29),
    .din_7_30(din_7_30_r2),
    .din_valid_7_30(din_valid_7_30_r2),
    .din_almost_full_7_30(din_almost_full_7_30),
    .din_7_31(din_7_31_r2),
    .din_valid_7_31(din_valid_7_31_r2),
    .din_almost_full_7_31(din_almost_full_7_31),
    .ruleID(out_data),
    .ruleID_valid(out_valid),
    .ruleID_last(out_last),
    .ruleID_almost_full(out_almost_full),
    .clk_status         (clk_status),
    .status_addr        (status_addr),
    .status_read        (status_read),
    .status_write       (status_write),
    .status_writedata   (status_writedata),
    .status_readdata    (status_readdata_back),
    .status_readdata_valid (status_readdata_valid_back)
);

endmodule //top